  // Interpreting sha_test.hex as an Intel formal HEX file.
  reg [7:0] rombuf[244:0];
  always @(posedge clk) begin
    if(rst) begin
      rombuf[0] = 8'h2;
      rombuf[1] = 8'h0;
      rombuf[2] = 8'h6;
      rombuf[3] = 8'h2;
      rombuf[4] = 8'h0;
      rombuf[5] = 8'h88;
      rombuf[6] = 8'h75;
      rombuf[7] = 8'h81;
      rombuf[8] = 8'h7;
      rombuf[9] = 8'h12;
      rombuf[10] = 8'h0;
      rombuf[11] = 8'hf1;
      rombuf[12] = 8'he5;
      rombuf[13] = 8'h82;
      rombuf[14] = 8'h60;
      rombuf[15] = 8'h3;
      rombuf[16] = 8'h2;
      rombuf[17] = 8'h0;
      rombuf[18] = 8'h3;
      rombuf[19] = 8'h79;
      rombuf[20] = 8'h0;
      rombuf[21] = 8'he9;
      rombuf[22] = 8'h44;
      rombuf[23] = 8'h0;
      rombuf[24] = 8'h60;
      rombuf[25] = 8'h1b;
      rombuf[26] = 8'h7a;
      rombuf[27] = 8'h0;
      rombuf[28] = 8'h90;
      rombuf[29] = 8'h0;
      rombuf[30] = 8'hf5;
      rombuf[31] = 8'h78;
      rombuf[32] = 8'h1;
      rombuf[33] = 8'h75;
      rombuf[34] = 8'ha0;
      rombuf[35] = 8'h0;
      rombuf[36] = 8'he4;
      rombuf[37] = 8'h93;
      rombuf[38] = 8'hf2;
      rombuf[39] = 8'ha3;
      rombuf[40] = 8'h8;
      rombuf[41] = 8'hb8;
      rombuf[42] = 8'h0;
      rombuf[43] = 8'h2;
      rombuf[44] = 8'h5;
      rombuf[45] = 8'ha0;
      rombuf[46] = 8'hd9;
      rombuf[47] = 8'hf4;
      rombuf[48] = 8'hda;
      rombuf[49] = 8'hf2;
      rombuf[50] = 8'h75;
      rombuf[51] = 8'ha0;
      rombuf[52] = 8'hff;
      rombuf[53] = 8'he4;
      rombuf[54] = 8'h78;
      rombuf[55] = 8'hff;
      rombuf[56] = 8'hf6;
      rombuf[57] = 8'hd8;
      rombuf[58] = 8'hfd;
      rombuf[59] = 8'h78;
      rombuf[60] = 8'h0;
      rombuf[61] = 8'he8;
      rombuf[62] = 8'h44;
      rombuf[63] = 8'h0;
      rombuf[64] = 8'h60;
      rombuf[65] = 8'ha;
      rombuf[66] = 8'h79;
      rombuf[67] = 8'h1;
      rombuf[68] = 8'h75;
      rombuf[69] = 8'ha0;
      rombuf[70] = 8'h0;
      rombuf[71] = 8'he4;
      rombuf[72] = 8'hf3;
      rombuf[73] = 8'h9;
      rombuf[74] = 8'hd8;
      rombuf[75] = 8'hfc;
      rombuf[76] = 8'h78;
      rombuf[77] = 8'h0;
      rombuf[78] = 8'he8;
      rombuf[79] = 8'h44;
      rombuf[80] = 8'h0;
      rombuf[81] = 8'h60;
      rombuf[82] = 8'hc;
      rombuf[83] = 8'h79;
      rombuf[84] = 8'h0;
      rombuf[85] = 8'h90;
      rombuf[86] = 8'h0;
      rombuf[87] = 8'h1;
      rombuf[88] = 8'he4;
      rombuf[89] = 8'hf0;
      rombuf[90] = 8'ha3;
      rombuf[91] = 8'hd8;
      rombuf[92] = 8'hfc;
      rombuf[93] = 8'hd9;
      rombuf[94] = 8'hfa;
      rombuf[95] = 8'h2;
      rombuf[96] = 8'h0;
      rombuf[97] = 8'h3;
      rombuf[98] = 8'h75;
      rombuf[99] = 8'hb0;
      rombuf[100] = 8'hde;
      rombuf[101] = 8'h75;
      rombuf[102] = 8'ha0;
      rombuf[103] = 8'hde;
      rombuf[104] = 8'h75;
      rombuf[105] = 8'h90;
      rombuf[106] = 8'hde;
      rombuf[107] = 8'h75;
      rombuf[108] = 8'h80;
      rombuf[109] = 8'hde;
      rombuf[110] = 8'h75;
      rombuf[111] = 8'hb0;
      rombuf[112] = 8'had;
      rombuf[113] = 8'h75;
      rombuf[114] = 8'ha0;
      rombuf[115] = 8'had;
      rombuf[116] = 8'h75;
      rombuf[117] = 8'h90;
      rombuf[118] = 8'had;
      rombuf[119] = 8'h75;
      rombuf[120] = 8'h80;
      rombuf[121] = 8'had;
      rombuf[122] = 8'h75;
      rombuf[123] = 8'hb0;
      rombuf[124] = 8'h0;
      rombuf[125] = 8'h75;
      rombuf[126] = 8'ha0;
      rombuf[127] = 8'h0;
      rombuf[128] = 8'h75;
      rombuf[129] = 8'h90;
      rombuf[130] = 8'h0;
      rombuf[131] = 8'h75;
      rombuf[132] = 8'h80;
      rombuf[133] = 8'h0;
      rombuf[134] = 8'h80;
      rombuf[135] = 8'hfe;
      rombuf[136] = 8'h7e;
      rombuf[137] = 8'h0;
      rombuf[138] = 8'h7f;
      rombuf[139] = 8'h0;
      rombuf[140] = 8'h8e;
      rombuf[141] = 8'h82;
      rombuf[142] = 8'h74;
      rombuf[143] = 8'he0;
      rombuf[144] = 8'h2f;
      rombuf[145] = 8'hf5;
      rombuf[146] = 8'h83;
      rombuf[147] = 8'h8e;
      rombuf[148] = 8'h5;
      rombuf[149] = 8'hed;
      rombuf[150] = 8'hf0;
      rombuf[151] = 8'he;
      rombuf[152] = 8'hbe;
      rombuf[153] = 8'h0;
      rombuf[154] = 8'h1;
      rombuf[155] = 8'hf;
      rombuf[156] = 8'hc3;
      rombuf[157] = 8'hee;
      rombuf[158] = 8'h94;
      rombuf[159] = 8'h20;
      rombuf[160] = 8'hef;
      rombuf[161] = 8'h64;
      rombuf[162] = 8'h80;
      rombuf[163] = 8'h94;
      rombuf[164] = 8'h80;
      rombuf[165] = 8'h40;
      rombuf[166] = 8'he5;
      rombuf[167] = 8'h90;
      rombuf[168] = 8'hfe;
      rombuf[169] = 8'h2;
      rombuf[170] = 8'h74;
      rombuf[171] = 8'h0;
      rombuf[172] = 8'hf0;
      rombuf[173] = 8'h74;
      rombuf[174] = 8'he0;
      rombuf[175] = 8'ha3;
      rombuf[176] = 8'hf0;
      rombuf[177] = 8'h90;
      rombuf[178] = 8'hfe;
      rombuf[179] = 8'h4;
      rombuf[180] = 8'h74;
      rombuf[181] = 8'h0;
      rombuf[182] = 8'hf0;
      rombuf[183] = 8'h74;
      rombuf[184] = 8'he1;
      rombuf[185] = 8'ha3;
      rombuf[186] = 8'hf0;
      rombuf[187] = 8'h90;
      rombuf[188] = 8'hfe;
      rombuf[189] = 8'h6;
      rombuf[190] = 8'h74;
      rombuf[191] = 8'h20;
      rombuf[192] = 8'hf0;
      rombuf[193] = 8'he4;
      rombuf[194] = 8'ha3;
      rombuf[195] = 8'hf0;
      rombuf[196] = 8'h90;
      rombuf[197] = 8'hfe;
      rombuf[198] = 8'h0;
      rombuf[199] = 8'h4;
      rombuf[200] = 8'hf0;
      rombuf[201] = 8'h90;
      rombuf[202] = 8'hfe;
      rombuf[203] = 8'h1;
      rombuf[204] = 8'he0;
      rombuf[205] = 8'hff;
      rombuf[206] = 8'h70;
      rombuf[207] = 8'hf9;
      rombuf[208] = 8'hfe;
      rombuf[209] = 8'hff;
      rombuf[210] = 8'h8e;
      rombuf[211] = 8'h90;
      rombuf[212] = 8'h8e;
      rombuf[213] = 8'h82;
      rombuf[214] = 8'h74;
      rombuf[215] = 8'he1;
      rombuf[216] = 8'h2f;
      rombuf[217] = 8'hf5;
      rombuf[218] = 8'h83;
      rombuf[219] = 8'he0;
      rombuf[220] = 8'hf5;
      rombuf[221] = 8'h80;
      rombuf[222] = 8'he;
      rombuf[223] = 8'hbe;
      rombuf[224] = 8'h0;
      rombuf[225] = 8'h1;
      rombuf[226] = 8'hf;
      rombuf[227] = 8'hc3;
      rombuf[228] = 8'hee;
      rombuf[229] = 8'h94;
      rombuf[230] = 8'h14;
      rombuf[231] = 8'hef;
      rombuf[232] = 8'h64;
      rombuf[233] = 8'h80;
      rombuf[234] = 8'h94;
      rombuf[235] = 8'h80;
      rombuf[236] = 8'h40;
      rombuf[237] = 8'he4;
      rombuf[238] = 8'h2;
      rombuf[239] = 8'h0;
      rombuf[240] = 8'h62;
      rombuf[241] = 8'h75;
      rombuf[242] = 8'h82;
      rombuf[243] = 8'h0;
      rombuf[244] = 8'h22;
    end
  end
  wire [15:0] addr0 = addr;
  wire [15:0] addr1 = addr+1;
  wire [15:0] addr2 = addr+2;
  wire [15:0] addr3 = addr+3;
  wire [7:0] data_o0 = (addr0 < 245) ? rombuf[addr0] : 8'hx;
  wire [7:0] data_o1 = (addr1 < 245) ? rombuf[addr1] : 8'hx;
  wire [7:0] data_o2 = (addr2 < 245) ? rombuf[addr2] : 8'hx;
  wire [7:0] data_o3 = (addr3 < 245) ? rombuf[addr3] : 8'hx;
  wire [31:0] data_out = {data_o3, data_o2, data_o1, data_o0};
