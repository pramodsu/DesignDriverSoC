
  reg [7:0] rombuf[64:0];
  always @(posedge clk) begin
    if(rst) begin
      rombuf[0] = 8'hx;
      rombuf[1] = 8'hx;
      rombuf[2] = 8'hx;
      rombuf[3] = 8'hx;
      rombuf[4] = 8'hx;
      rombuf[5] = 8'hx;
      rombuf[6] = 8'hx;
      rombuf[7] = 8'hx;
      rombuf[8] = 8'hx;
      rombuf[9] = 8'hx;
      rombuf[10] = 8'hx;
      rombuf[11] = 8'hx;
      rombuf[12] = 8'hx;
      rombuf[13] = 8'hx;
      rombuf[14] = 8'hx;
      rombuf[15] = 8'hx;
      rombuf[16] = 8'hx;
      rombuf[17] = 8'hx;
      rombuf[18] = 8'hx;
      rombuf[19] = 8'hx;
      rombuf[20] = 8'hx;
      rombuf[21] = 8'hx;
      rombuf[22] = 8'hx;
      rombuf[23] = 8'hx;
      rombuf[24] = 8'hx;
      rombuf[25] = 8'hx;
      rombuf[26] = 8'hx;
      rombuf[27] = 8'hx;
      rombuf[28] = 8'hx;
      rombuf[29] = 8'hx;
      rombuf[30] = 8'hx;
      rombuf[31] = 8'hx;
      rombuf[32] = 8'hx;
      rombuf[33] = 8'hx;
      rombuf[34] = 8'hx;
      rombuf[35] = 8'hx;
      rombuf[36] = 8'hx;
      rombuf[37] = 8'hx;
      rombuf[38] = 8'hx;
      rombuf[39] = 8'hx;
      rombuf[40] = 8'hx;
      rombuf[41] = 8'hx;
      rombuf[42] = 8'hx;
      rombuf[43] = 8'hx;
      rombuf[44] = 8'hx;
      rombuf[45] = 8'hx;
      rombuf[46] = 8'hx;
      rombuf[47] = 8'hx;
      rombuf[48] = 8'hx;
      rombuf[49] = 8'hx;
      rombuf[50] = 8'hx;
      rombuf[51] = 8'hx;
      rombuf[52] = 8'hx;
      rombuf[53] = 8'hx;
      rombuf[54] = 8'hx;
      rombuf[55] = 8'hx;
      rombuf[56] = 8'hx;
      rombuf[57] = 8'hx;
      rombuf[58] = 8'hx;
      rombuf[59] = 8'hx;
      rombuf[60] = 8'hx;
      rombuf[61] = 8'hx;
      rombuf[62] = 8'hx;
      rombuf[63] = 8'hx;
    end
  end
  wire [15:0] addr0 = addr;
  wire [15:0] addr1 = addr+1;
  wire [15:0] addr2 = addr+2;
  wire [15:0] addr3 = addr+3;
  wire [7:0] data_o0 = (addr0 < 64) ? rombuf[addr0] : 8'hx;
  wire [7:0] data_o1 = (addr1 < 64) ? rombuf[addr1] : 8'hx;
  wire [7:0] data_o2 = (addr2 < 64) ? rombuf[addr2] : 8'hx;
  wire [7:0] data_o3 = (addr3 < 64) ? rombuf[addr3] : 8'hx;
  wire [31:0] data_out = {data_o3, data_o2, data_o1, data_o0};
