module xm8051_golden_model(
  clk,
  rst,
  step,
  RD_xram_0_ADDR,
  RD_xram_1_ADDR,
  RD_xram_2_ADDR,
  RD_xram_3_ADDR,
  RD_xram_4_ADDR,
  RD_xram_5_ADDR,
  RD_xram_6_ADDR,
  RD_xram_7_ADDR,
  RD_xram_8_ADDR,
  RD_xram_9_ADDR,
  RD_xram_10_ADDR,
  RD_xram_11_ADDR,
  RD_xram_12_ADDR,
  RD_xram_13_ADDR,
  RD_xram_14_ADDR,
  RD_xram_15_ADDR,
  RD_xram_16_ADDR,
  RD_xram_17_ADDR,
  RD_xram_18_ADDR,
  RD_xram_19_ADDR,
  RD_xram_20_ADDR,
  RD_xram_21_ADDR,
  RD_xram_22_ADDR,
  RD_xram_23_ADDR,
  RD_xram_24_ADDR,
  RD_xram_25_ADDR,
  RD_xram_26_ADDR,
  RD_xram_27_ADDR,
  RD_xram_28_ADDR,
  RD_xram_29_ADDR,
  RD_xram_30_ADDR,
  RD_xram_31_ADDR,
  RD_xram_32_ADDR,
  RD_xram_33_ADDR,
  RD_xram_34_ADDR,
  RD_xram_35_ADDR,
  RD_xram_36_ADDR,
  RD_xram_37_ADDR,
  RD_xram_38_ADDR,
  RD_xram_39_ADDR,
  RD_xram_40_ADDR,
  RD_xram_41_ADDR,
  RD_xram_42_ADDR,
  RD_xram_43_ADDR,
  RD_xram_44_ADDR,
  RD_xram_45_ADDR,
  RD_xram_46_ADDR,
  RD_xram_47_ADDR,
  RD_xram_48_ADDR,
  RD_xram_49_ADDR,
  RD_xram_50_ADDR,
  RD_xram_51_ADDR,
  RD_xram_52_ADDR,
  RD_xram_53_ADDR,
  RD_xram_54_ADDR,
  RD_xram_55_ADDR,
  RD_xram_56_ADDR,
  RD_xram_57_ADDR,
  RD_xram_58_ADDR,
  RD_xram_59_ADDR,
  RD_xram_60_ADDR,
  RD_xram_61_ADDR,
  RD_xram_62_ADDR,
  RD_xram_63_ADDR,
  RD_xram_64_ADDR,
  RD_xram_65_ADDR,
  RD_xram_66_ADDR,
  RD_xram_67_ADDR,
  RD_xram_68_ADDR,
  RD_xram_69_ADDR,
  RD_xram_70_ADDR,
  RD_xram_71_ADDR,
  RD_xram_72_ADDR,
  RD_xram_73_ADDR,
  RD_xram_74_ADDR,
  RD_xram_75_ADDR,
  RD_xram_76_ADDR,
  RD_xram_77_ADDR,
  RD_xram_78_ADDR,
  RD_xram_79_ADDR,
  RD_xram_80_ADDR,
  sha_read_data,
  sha_read_data_next,
  aes_read_data,
  aes_read_data_next,
  sha_rdaddr,
  sha_rdaddr_next,
  aes_addr,
  aes_addr_next,
  aes_ctr,
  aes_ctr_next,
  aes_bytes_processed,
  aes_bytes_processed_next,
  sha_len,
  sha_len_next,
  aes_key1,
  aes_key1_next,
  aes_key0,
  aes_key0_next,
  aes_len,
  aes_len_next,
  sha_bytes_processed,
  sha_bytes_processed_next,
  sha_wraddr,
  sha_wraddr_next,
  dataout,
  dataout_next,
  WR_XRAM_ADDR,
  WR_XRAM_ADDR_next,
  WR_XRAM_EN,
  WR_XRAM_EN_next,
  aes_state,
  aes_state_next,
  aes_enc_data,
  aes_enc_data_next,
  sha_state,
  sha_state_next,
  sha_digest,
  sha_digest_next,
  op,
  addrin,
  datain,
  input_sha_func_0,
  input_sha_func_1,
  input_sha_func_2,
  input_sha_func_3,
  input_sha_func_4,
  input_sha_func_5,
  input_aes_func_6,
  input_aes_func_7,
  input_sha_func_8,
  input_sha_func_9,
  input_sha_func_10,
  input_sha_func_11,
  input_sha_func_12,
  input_sha_func_13,
  input_sha_func_14,
  input_sha_func_15,
  input_sha_func_16,
  input_sha_func_17,
  input_sha_func_18,
  input_sha_func_19,
  input_sha_func_20,
  input_sha_func_21,
  input_sha_func_22,
  input_aes_func_23,
  input_aes_func_24,
  input_sha_func_25,
  input_sha_func_26,
  input_sha_func_27,
  input_sha_func_28,
  input_sha_func_29,
  input_sha_func_30,
  input_sha_func_31,
  input_sha_func_32,
  input_sha_func_33,
  input_sha_func_34,
  input_sha_func_35,
  input_sha_func_36,
  input_aes_func_37,
  input_aes_func_38,
  input_sha_func_39,
  input_sha_func_40,
  input_sha_func_41,
  input_sha_func_42,
  input_sha_func_43,
  input_sha_func_44,
  input_sha_func_45,
  input_sha_func_46,
  input_sha_func_47,
  input_sha_func_48,
  input_sha_func_49,
  input_sha_func_50,
  input_aes_func_51,
  input_aes_func_52,
  input_sha_func_53,
  input_sha_func_54,
  input_sha_func_55,
  RD_xram_0,
  RD_xram_1,
  RD_xram_2,
  RD_xram_3,
  RD_xram_4,
  RD_xram_5,
  RD_xram_6,
  RD_xram_7,
  RD_xram_8,
  RD_xram_9,
  RD_xram_10,
  RD_xram_11,
  RD_xram_12,
  RD_xram_13,
  RD_xram_14,
  RD_xram_15,
  RD_xram_16,
  RD_xram_17,
  RD_xram_18,
  RD_xram_19,
  RD_xram_20,
  RD_xram_21,
  RD_xram_22,
  RD_xram_23,
  RD_xram_24,
  RD_xram_25,
  RD_xram_26,
  RD_xram_27,
  RD_xram_28,
  RD_xram_29,
  RD_xram_30,
  RD_xram_31,
  RD_xram_32,
  RD_xram_33,
  RD_xram_34,
  RD_xram_35,
  RD_xram_36,
  RD_xram_37,
  RD_xram_38,
  RD_xram_39,
  RD_xram_40,
  RD_xram_41,
  RD_xram_42,
  RD_xram_43,
  RD_xram_44,
  RD_xram_45,
  RD_xram_46,
  RD_xram_47,
  RD_xram_48,
  RD_xram_49,
  RD_xram_50,
  RD_xram_51,
  RD_xram_52,
  RD_xram_53,
  RD_xram_54,
  RD_xram_55,
  RD_xram_56,
  RD_xram_57,
  RD_xram_58,
  RD_xram_59,
  RD_xram_60,
  RD_xram_61,
  RD_xram_62,
  RD_xram_63,
  RD_xram_64,
  RD_xram_65,
  RD_xram_66,
  RD_xram_67,
  RD_xram_68,
  RD_xram_69,
  RD_xram_70,
  RD_xram_71,
  RD_xram_72,
  RD_xram_73,
  RD_xram_74,
  RD_xram_75,
  RD_xram_76,
  RD_xram_77,
  RD_xram_78,
  RD_xram_79,
  RD_xram_80,
  nondet_memwrite_choice_0,
  nondet_memwrite_choice_1,
  nondet_memwrite_choice_2,
  nondet_memwrite_choice_3,
  nondet_memwrite_choice_4,
  nondet_memwrite_choice_5,
  nondet_memwrite_choice_6,
  nondet_memwrite_choice_7,
  nondet_memwrite_choice_8,
  nondet_memwrite_choice_9,
  nondet_memwrite_choice_10,
  nondet_memwrite_choice_11,
  nondet_memwrite_choice_12,
  nondet_memwrite_choice_13,
  nondet_memwrite_choice_14,
  nondet_memwrite_choice_15,
  nondet_memwrite_choice_16,
  nondet_memwrite_choice_17,
  nondet_memwrite_choice_18,
  nondet_memwrite_choice_19,
  nondet_memwrite_choice_20,
  nondet_memwrite_choice_21,
  nondet_memwrite_choice_22,
  nondet_memwrite_choice_23,
  nondet_memwrite_choice_24,
  nondet_memwrite_choice_25,
  nondet_memwrite_choice_26,
  nondet_memwrite_choice_27,
  nondet_memwrite_choice_28,
  nondet_memwrite_choice_29,
  nondet_memwrite_choice_30,
  nondet_memwrite_choice_31,
  nondet_memwrite_choice_32,
  nondet_memwrite_choice_33,
  nondet_memwrite_choice_34,
  nondet_memwrite_choice_35,
  nondet_memwrite_choice_36,
  nondet_memwrite_choice_37,
  nondet_memwrite_choice_38,
  nondet_memwrite_choice_39,
  nondet_memwrite_choice_40,
  nondet_memwrite_choice_41,
  nondet_memwrite_choice_42,
  nondet_memwrite_choice_43,
  nondet_memwrite_choice_44,
  nondet_memwrite_choice_45,
  nondet_memwrite_choice_46,
  nondet_memwrite_choice_47,
  nondet_memwrite_choice_48,
  nondet_memwrite_choice_49,
  nondet_memwrite_choice_50,
  nondet_memwrite_choice_51,
  nondet_memwrite_choice_52,
  nondet_memwrite_choice_53,
  nondet_memwrite_choice_54,
  nondet_memwrite_choice_55,
  nondet_memwrite_choice_56,
  nondet_memwrite_choice_57,
  nondet_memwrite_choice_58,
  nondet_memwrite_choice_59,
  nondet_memwrite_choice_60,
  nondet_memwrite_choice_61,
  nondet_memwrite_choice_62,
  nondet_memwrite_choice_63,
  nondet_memwrite_choice_64,
  nondet_memwrite_choice_65,
  nondet_memwrite_choice_66,
  nondet_memwrite_choice_67,
  nondet_memwrite_choice_68,
  nondet_memwrite_choice_69,
  nondet_memwrite_choice_70,
  nondet_memwrite_choice_71,
  nondet_memwrite_choice_72,
  nondet_memwrite_choice_73,
  nondet_memwrite_choice_74,
  nondet_memwrite_choice_75,
  nondet_memwrite_choice_76,
  nondet_memwrite_choice_77,
  nondet_memwrite_choice_78,
  nondet_memwrite_choice_79,
  nondet_memwrite_choice_80,
  nondet_memwrite_choice_81,
  nondet_memwrite_choice_82,
  nondet_memwrite_choice_83,
  nondet_memwrite_choice_84,
  nondet_memwrite_choice_85,
  nondet_memwrite_choice_86,
  nondet_memwrite_choice_87,
  nondet_memwrite_choice_88,
  nondet_memwrite_choice_89,
  nondet_memwrite_choice_90,
  nondet_memwrite_choice_91,
  nondet_memwrite_choice_92,
  nondet_memwrite_choice_93,
  nondet_memwrite_choice_94,
  nondet_memwrite_choice_95,
  nondet_memwrite_choice_96,
  nondet_memwrite_choice_97,
  nondet_memwrite_choice_98,
  nondet_memwrite_choice_99,
  nondet_memwrite_choice_100,
  nondet_memwrite_choice_101,
  nondet_memwrite_choice_102,
  nondet_memwrite_choice_103,
  nondet_memwrite_choice_104,
  nondet_memwrite_choice_105,
  nondet_memwrite_choice_106,
  nondet_memwrite_choice_107,
  nondet_memwrite_choice_108,
  nondet_memwrite_choice_109,
  nondet_memwrite_choice_110,
  nondet_memwrite_choice_111,
  nondet_memwrite_choice_112,
  nondet_memwrite_choice_113,
  nondet_memwrite_choice_114,
  nondet_memwrite_choice_115,
  nondet_memwrite_choice_116,
  nondet_memwrite_choice_117,
  nondet_memwrite_choice_118,
  nondet_memwrite_choice_119
);
output [15:0] RD_xram_0_ADDR;
output [15:0] RD_xram_1_ADDR;
output [15:0] RD_xram_2_ADDR;
output [15:0] RD_xram_3_ADDR;
output [15:0] RD_xram_4_ADDR;
output [15:0] RD_xram_5_ADDR;
output [15:0] RD_xram_6_ADDR;
output [15:0] RD_xram_7_ADDR;
output [15:0] RD_xram_8_ADDR;
output [15:0] RD_xram_9_ADDR;
output [15:0] RD_xram_10_ADDR;
output [15:0] RD_xram_11_ADDR;
output [15:0] RD_xram_12_ADDR;
output [15:0] RD_xram_13_ADDR;
output [15:0] RD_xram_14_ADDR;
output [15:0] RD_xram_15_ADDR;
output [15:0] RD_xram_16_ADDR;
output [15:0] RD_xram_17_ADDR;
output [15:0] RD_xram_18_ADDR;
output [15:0] RD_xram_19_ADDR;
output [15:0] RD_xram_20_ADDR;
output [15:0] RD_xram_21_ADDR;
output [15:0] RD_xram_22_ADDR;
output [15:0] RD_xram_23_ADDR;
output [15:0] RD_xram_24_ADDR;
output [15:0] RD_xram_25_ADDR;
output [15:0] RD_xram_26_ADDR;
output [15:0] RD_xram_27_ADDR;
output [15:0] RD_xram_28_ADDR;
output [15:0] RD_xram_29_ADDR;
output [15:0] RD_xram_30_ADDR;
output [15:0] RD_xram_31_ADDR;
output [15:0] RD_xram_32_ADDR;
output [15:0] RD_xram_33_ADDR;
output [15:0] RD_xram_34_ADDR;
output [15:0] RD_xram_35_ADDR;
output [15:0] RD_xram_36_ADDR;
output [15:0] RD_xram_37_ADDR;
output [15:0] RD_xram_38_ADDR;
output [15:0] RD_xram_39_ADDR;
output [15:0] RD_xram_40_ADDR;
output [15:0] RD_xram_41_ADDR;
output [15:0] RD_xram_42_ADDR;
output [15:0] RD_xram_43_ADDR;
output [15:0] RD_xram_44_ADDR;
output [15:0] RD_xram_45_ADDR;
output [15:0] RD_xram_46_ADDR;
output [15:0] RD_xram_47_ADDR;
output [15:0] RD_xram_48_ADDR;
output [15:0] RD_xram_49_ADDR;
output [15:0] RD_xram_50_ADDR;
output [15:0] RD_xram_51_ADDR;
output [15:0] RD_xram_52_ADDR;
output [15:0] RD_xram_53_ADDR;
output [15:0] RD_xram_54_ADDR;
output [15:0] RD_xram_55_ADDR;
output [15:0] RD_xram_56_ADDR;
output [15:0] RD_xram_57_ADDR;
output [15:0] RD_xram_58_ADDR;
output [15:0] RD_xram_59_ADDR;
output [15:0] RD_xram_60_ADDR;
output [15:0] RD_xram_61_ADDR;
output [15:0] RD_xram_62_ADDR;
output [15:0] RD_xram_63_ADDR;
output [15:0] RD_xram_64_ADDR;
output [15:0] RD_xram_65_ADDR;
output [15:0] RD_xram_66_ADDR;
output [15:0] RD_xram_67_ADDR;
output [15:0] RD_xram_68_ADDR;
output [15:0] RD_xram_69_ADDR;
output [15:0] RD_xram_70_ADDR;
output [15:0] RD_xram_71_ADDR;
output [15:0] RD_xram_72_ADDR;
output [15:0] RD_xram_73_ADDR;
output [15:0] RD_xram_74_ADDR;
output [15:0] RD_xram_75_ADDR;
output [15:0] RD_xram_76_ADDR;
output [15:0] RD_xram_77_ADDR;
output [15:0] RD_xram_78_ADDR;
output [15:0] RD_xram_79_ADDR;
output [15:0] RD_xram_80_ADDR;
output [511:0] sha_read_data;
output [511:0] sha_read_data_next;
output [127:0] aes_read_data;
output [127:0] aes_read_data_next;
output [15:0] sha_rdaddr;
output [15:0] sha_rdaddr_next;
output [15:0] aes_addr;
output [15:0] aes_addr_next;
output [127:0] aes_ctr;
output [127:0] aes_ctr_next;
output [15:0] aes_bytes_processed;
output [15:0] aes_bytes_processed_next;
output [15:0] sha_len;
output [15:0] sha_len_next;
output [127:0] aes_key1;
output [127:0] aes_key1_next;
output [127:0] aes_key0;
output [127:0] aes_key0_next;
output [15:0] aes_len;
output [15:0] aes_len_next;
output [15:0] sha_bytes_processed;
output [15:0] sha_bytes_processed_next;
output [15:0] sha_wraddr;
output [15:0] sha_wraddr_next;
output [7:0] dataout;
output [7:0] dataout_next;
output [15:0] WR_XRAM_ADDR;
output [15:0] WR_XRAM_ADDR_next;
output WR_XRAM_EN;
output WR_XRAM_EN_next;
output [7:0] aes_state;
output [7:0] aes_state_next;
output [127:0] aes_enc_data;
output [127:0] aes_enc_data_next;
output [7:0] sha_state;
output [7:0] sha_state_next;
output [159:0] sha_digest;
output [159:0] sha_digest_next;

input clk, rst, step;
input [3:0] op;
input [15:0] addrin;
input [7:0] datain;
input [63:0] input_sha_func_0;
input [63:0] input_sha_func_1;
input [31:0] input_sha_func_2;
input [63:0] input_sha_func_3;
input [63:0] input_sha_func_4;
input [31:0] input_sha_func_5;
input [63:0] input_aes_func_6;
input [63:0] input_aes_func_7;
input [63:0] input_sha_func_8;
input [63:0] input_sha_func_9;
input [31:0] input_sha_func_10;
input [63:0] input_sha_func_11;
input [63:0] input_sha_func_12;
input [31:0] input_sha_func_13;
input [63:0] input_sha_func_14;
input [63:0] input_sha_func_15;
input [31:0] input_sha_func_16;
input [63:0] input_sha_func_17;
input [63:0] input_sha_func_18;
input [31:0] input_sha_func_19;
input [63:0] input_sha_func_20;
input [63:0] input_sha_func_21;
input [31:0] input_sha_func_22;
input [63:0] input_aes_func_23;
input [63:0] input_aes_func_24;
input [63:0] input_sha_func_25;
input [63:0] input_sha_func_26;
input [31:0] input_sha_func_27;
input [63:0] input_sha_func_28;
input [63:0] input_sha_func_29;
input [31:0] input_sha_func_30;
input [63:0] input_sha_func_31;
input [63:0] input_sha_func_32;
input [31:0] input_sha_func_33;
input [63:0] input_sha_func_34;
input [63:0] input_sha_func_35;
input [31:0] input_sha_func_36;
input [63:0] input_aes_func_37;
input [63:0] input_aes_func_38;
input [63:0] input_sha_func_39;
input [63:0] input_sha_func_40;
input [31:0] input_sha_func_41;
input [63:0] input_sha_func_42;
input [63:0] input_sha_func_43;
input [31:0] input_sha_func_44;
input [63:0] input_sha_func_45;
input [63:0] input_sha_func_46;
input [31:0] input_sha_func_47;
input [63:0] input_sha_func_48;
input [63:0] input_sha_func_49;
input [31:0] input_sha_func_50;
input [63:0] input_aes_func_51;
input [63:0] input_aes_func_52;
input [63:0] input_sha_func_53;
input [63:0] input_sha_func_54;
input [31:0] input_sha_func_55;
input [7:0] RD_xram_0;
input [7:0] RD_xram_1;
input [7:0] RD_xram_2;
input [7:0] RD_xram_3;
input [7:0] RD_xram_4;
input [7:0] RD_xram_5;
input [7:0] RD_xram_6;
input [7:0] RD_xram_7;
input [7:0] RD_xram_8;
input [7:0] RD_xram_9;
input [7:0] RD_xram_10;
input [7:0] RD_xram_11;
input [7:0] RD_xram_12;
input [7:0] RD_xram_13;
input [7:0] RD_xram_14;
input [7:0] RD_xram_15;
input [7:0] RD_xram_16;
input [7:0] RD_xram_17;
input [7:0] RD_xram_18;
input [7:0] RD_xram_19;
input [7:0] RD_xram_20;
input [7:0] RD_xram_21;
input [7:0] RD_xram_22;
input [7:0] RD_xram_23;
input [7:0] RD_xram_24;
input [7:0] RD_xram_25;
input [7:0] RD_xram_26;
input [7:0] RD_xram_27;
input [7:0] RD_xram_28;
input [7:0] RD_xram_29;
input [7:0] RD_xram_30;
input [7:0] RD_xram_31;
input [7:0] RD_xram_32;
input [7:0] RD_xram_33;
input [7:0] RD_xram_34;
input [7:0] RD_xram_35;
input [7:0] RD_xram_36;
input [7:0] RD_xram_37;
input [7:0] RD_xram_38;
input [7:0] RD_xram_39;
input [7:0] RD_xram_40;
input [7:0] RD_xram_41;
input [7:0] RD_xram_42;
input [7:0] RD_xram_43;
input [7:0] RD_xram_44;
input [7:0] RD_xram_45;
input [7:0] RD_xram_46;
input [7:0] RD_xram_47;
input [7:0] RD_xram_48;
input [7:0] RD_xram_49;
input [7:0] RD_xram_50;
input [7:0] RD_xram_51;
input [7:0] RD_xram_52;
input [7:0] RD_xram_53;
input [7:0] RD_xram_54;
input [7:0] RD_xram_55;
input [7:0] RD_xram_56;
input [7:0] RD_xram_57;
input [7:0] RD_xram_58;
input [7:0] RD_xram_59;
input [7:0] RD_xram_60;
input [7:0] RD_xram_61;
input [7:0] RD_xram_62;
input [7:0] RD_xram_63;
input [7:0] RD_xram_64;
input [7:0] RD_xram_65;
input [7:0] RD_xram_66;
input [7:0] RD_xram_67;
input [7:0] RD_xram_68;
input [7:0] RD_xram_69;
input [7:0] RD_xram_70;
input [7:0] RD_xram_71;
input [7:0] RD_xram_72;
input [7:0] RD_xram_73;
input [7:0] RD_xram_74;
input [7:0] RD_xram_75;
input [7:0] RD_xram_76;
input [7:0] RD_xram_77;
input [7:0] RD_xram_78;
input [7:0] RD_xram_79;
input [7:0] RD_xram_80;
input nondet_memwrite_choice_0;
input nondet_memwrite_choice_1;
input nondet_memwrite_choice_2;
input nondet_memwrite_choice_3;
input nondet_memwrite_choice_4;
input nondet_memwrite_choice_5;
input nondet_memwrite_choice_6;
input nondet_memwrite_choice_7;
input nondet_memwrite_choice_8;
input nondet_memwrite_choice_9;
input nondet_memwrite_choice_10;
input nondet_memwrite_choice_11;
input nondet_memwrite_choice_12;
input nondet_memwrite_choice_13;
input nondet_memwrite_choice_14;
input nondet_memwrite_choice_15;
input nondet_memwrite_choice_16;
input nondet_memwrite_choice_17;
input nondet_memwrite_choice_18;
input nondet_memwrite_choice_19;
input nondet_memwrite_choice_20;
input nondet_memwrite_choice_21;
input nondet_memwrite_choice_22;
input nondet_memwrite_choice_23;
input nondet_memwrite_choice_24;
input nondet_memwrite_choice_25;
input nondet_memwrite_choice_26;
input nondet_memwrite_choice_27;
input nondet_memwrite_choice_28;
input nondet_memwrite_choice_29;
input nondet_memwrite_choice_30;
input nondet_memwrite_choice_31;
input nondet_memwrite_choice_32;
input nondet_memwrite_choice_33;
input nondet_memwrite_choice_34;
input nondet_memwrite_choice_35;
input nondet_memwrite_choice_36;
input nondet_memwrite_choice_37;
input nondet_memwrite_choice_38;
input nondet_memwrite_choice_39;
input nondet_memwrite_choice_40;
input nondet_memwrite_choice_41;
input nondet_memwrite_choice_42;
input nondet_memwrite_choice_43;
input nondet_memwrite_choice_44;
input nondet_memwrite_choice_45;
input nondet_memwrite_choice_46;
input nondet_memwrite_choice_47;
input nondet_memwrite_choice_48;
input nondet_memwrite_choice_49;
input nondet_memwrite_choice_50;
input nondet_memwrite_choice_51;
input nondet_memwrite_choice_52;
input nondet_memwrite_choice_53;
input nondet_memwrite_choice_54;
input nondet_memwrite_choice_55;
input nondet_memwrite_choice_56;
input nondet_memwrite_choice_57;
input nondet_memwrite_choice_58;
input nondet_memwrite_choice_59;
input nondet_memwrite_choice_60;
input nondet_memwrite_choice_61;
input nondet_memwrite_choice_62;
input nondet_memwrite_choice_63;
input nondet_memwrite_choice_64;
input nondet_memwrite_choice_65;
input nondet_memwrite_choice_66;
input nondet_memwrite_choice_67;
input nondet_memwrite_choice_68;
input nondet_memwrite_choice_69;
input nondet_memwrite_choice_70;
input nondet_memwrite_choice_71;
input nondet_memwrite_choice_72;
input nondet_memwrite_choice_73;
input nondet_memwrite_choice_74;
input nondet_memwrite_choice_75;
input nondet_memwrite_choice_76;
input nondet_memwrite_choice_77;
input nondet_memwrite_choice_78;
input nondet_memwrite_choice_79;
input nondet_memwrite_choice_80;
input nondet_memwrite_choice_81;
input nondet_memwrite_choice_82;
input nondet_memwrite_choice_83;
input nondet_memwrite_choice_84;
input nondet_memwrite_choice_85;
input nondet_memwrite_choice_86;
input nondet_memwrite_choice_87;
input nondet_memwrite_choice_88;
input nondet_memwrite_choice_89;
input nondet_memwrite_choice_90;
input nondet_memwrite_choice_91;
input nondet_memwrite_choice_92;
input nondet_memwrite_choice_93;
input nondet_memwrite_choice_94;
input nondet_memwrite_choice_95;
input nondet_memwrite_choice_96;
input nondet_memwrite_choice_97;
input nondet_memwrite_choice_98;
input nondet_memwrite_choice_99;
input nondet_memwrite_choice_100;
input nondet_memwrite_choice_101;
input nondet_memwrite_choice_102;
input nondet_memwrite_choice_103;
input nondet_memwrite_choice_104;
input nondet_memwrite_choice_105;
input nondet_memwrite_choice_106;
input nondet_memwrite_choice_107;
input nondet_memwrite_choice_108;
input nondet_memwrite_choice_109;
input nondet_memwrite_choice_110;
input nondet_memwrite_choice_111;
input nondet_memwrite_choice_112;
input nondet_memwrite_choice_113;
input nondet_memwrite_choice_114;
input nondet_memwrite_choice_115;
input nondet_memwrite_choice_116;
input nondet_memwrite_choice_117;
input nondet_memwrite_choice_118;
input nondet_memwrite_choice_119;

reg [15:0] WR_XRAM_ADDR;
reg WR_XRAM_EN;
reg [15:0] aes_addr;
reg [15:0] aes_bytes_processed;
reg [127:0] aes_ctr;
reg [127:0] aes_enc_data;
reg [127:0] aes_key0;
reg [127:0] aes_key1;
reg [15:0] aes_len;
reg [127:0] aes_read_data;
reg [7:0] aes_state;
reg [7:0] dataout;
reg [15:0] sha_bytes_processed;
reg [159:0] sha_digest;
reg [15:0] sha_len;
reg [15:0] sha_rdaddr;
reg [511:0] sha_read_data;
reg [7:0] sha_state;
reg [15:0] sha_wraddr;

wire [7:0] RD_xram_0;
wire [15:0] RD_xram_0_ADDR;
wire [7:0] RD_xram_1;
wire [7:0] RD_xram_10;
wire [15:0] RD_xram_10_ADDR;
wire [7:0] RD_xram_11;
wire [15:0] RD_xram_11_ADDR;
wire [7:0] RD_xram_12;
wire [15:0] RD_xram_12_ADDR;
wire [7:0] RD_xram_13;
wire [15:0] RD_xram_13_ADDR;
wire [7:0] RD_xram_14;
wire [15:0] RD_xram_14_ADDR;
wire [7:0] RD_xram_15;
wire [15:0] RD_xram_15_ADDR;
wire [7:0] RD_xram_16;
wire [15:0] RD_xram_16_ADDR;
wire [7:0] RD_xram_17;
wire [15:0] RD_xram_17_ADDR;
wire [7:0] RD_xram_18;
wire [15:0] RD_xram_18_ADDR;
wire [7:0] RD_xram_19;
wire [15:0] RD_xram_19_ADDR;
wire [15:0] RD_xram_1_ADDR;
wire [7:0] RD_xram_2;
wire [7:0] RD_xram_20;
wire [15:0] RD_xram_20_ADDR;
wire [7:0] RD_xram_21;
wire [15:0] RD_xram_21_ADDR;
wire [7:0] RD_xram_22;
wire [15:0] RD_xram_22_ADDR;
wire [7:0] RD_xram_23;
wire [15:0] RD_xram_23_ADDR;
wire [7:0] RD_xram_24;
wire [15:0] RD_xram_24_ADDR;
wire [7:0] RD_xram_25;
wire [15:0] RD_xram_25_ADDR;
wire [7:0] RD_xram_26;
wire [15:0] RD_xram_26_ADDR;
wire [7:0] RD_xram_27;
wire [15:0] RD_xram_27_ADDR;
wire [7:0] RD_xram_28;
wire [15:0] RD_xram_28_ADDR;
wire [7:0] RD_xram_29;
wire [15:0] RD_xram_29_ADDR;
wire [15:0] RD_xram_2_ADDR;
wire [7:0] RD_xram_3;
wire [7:0] RD_xram_30;
wire [15:0] RD_xram_30_ADDR;
wire [7:0] RD_xram_31;
wire [15:0] RD_xram_31_ADDR;
wire [7:0] RD_xram_32;
wire [15:0] RD_xram_32_ADDR;
wire [7:0] RD_xram_33;
wire [15:0] RD_xram_33_ADDR;
wire [7:0] RD_xram_34;
wire [15:0] RD_xram_34_ADDR;
wire [7:0] RD_xram_35;
wire [15:0] RD_xram_35_ADDR;
wire [7:0] RD_xram_36;
wire [15:0] RD_xram_36_ADDR;
wire [7:0] RD_xram_37;
wire [15:0] RD_xram_37_ADDR;
wire [7:0] RD_xram_38;
wire [15:0] RD_xram_38_ADDR;
wire [7:0] RD_xram_39;
wire [15:0] RD_xram_39_ADDR;
wire [15:0] RD_xram_3_ADDR;
wire [7:0] RD_xram_4;
wire [7:0] RD_xram_40;
wire [15:0] RD_xram_40_ADDR;
wire [7:0] RD_xram_41;
wire [15:0] RD_xram_41_ADDR;
wire [7:0] RD_xram_42;
wire [15:0] RD_xram_42_ADDR;
wire [7:0] RD_xram_43;
wire [15:0] RD_xram_43_ADDR;
wire [7:0] RD_xram_44;
wire [15:0] RD_xram_44_ADDR;
wire [7:0] RD_xram_45;
wire [15:0] RD_xram_45_ADDR;
wire [7:0] RD_xram_46;
wire [15:0] RD_xram_46_ADDR;
wire [7:0] RD_xram_47;
wire [15:0] RD_xram_47_ADDR;
wire [7:0] RD_xram_48;
wire [15:0] RD_xram_48_ADDR;
wire [7:0] RD_xram_49;
wire [15:0] RD_xram_49_ADDR;
wire [15:0] RD_xram_4_ADDR;
wire [7:0] RD_xram_5;
wire [7:0] RD_xram_50;
wire [15:0] RD_xram_50_ADDR;
wire [7:0] RD_xram_51;
wire [15:0] RD_xram_51_ADDR;
wire [7:0] RD_xram_52;
wire [15:0] RD_xram_52_ADDR;
wire [7:0] RD_xram_53;
wire [15:0] RD_xram_53_ADDR;
wire [7:0] RD_xram_54;
wire [15:0] RD_xram_54_ADDR;
wire [7:0] RD_xram_55;
wire [15:0] RD_xram_55_ADDR;
wire [7:0] RD_xram_56;
wire [15:0] RD_xram_56_ADDR;
wire [7:0] RD_xram_57;
wire [15:0] RD_xram_57_ADDR;
wire [7:0] RD_xram_58;
wire [15:0] RD_xram_58_ADDR;
wire [7:0] RD_xram_59;
wire [15:0] RD_xram_59_ADDR;
wire [15:0] RD_xram_5_ADDR;
wire [7:0] RD_xram_6;
wire [7:0] RD_xram_60;
wire [15:0] RD_xram_60_ADDR;
wire [7:0] RD_xram_61;
wire [15:0] RD_xram_61_ADDR;
wire [7:0] RD_xram_62;
wire [15:0] RD_xram_62_ADDR;
wire [7:0] RD_xram_63;
wire [15:0] RD_xram_63_ADDR;
wire [7:0] RD_xram_64;
wire [15:0] RD_xram_64_ADDR;
wire [7:0] RD_xram_65;
wire [15:0] RD_xram_65_ADDR;
wire [7:0] RD_xram_66;
wire [15:0] RD_xram_66_ADDR;
wire [7:0] RD_xram_67;
wire [15:0] RD_xram_67_ADDR;
wire [7:0] RD_xram_68;
wire [15:0] RD_xram_68_ADDR;
wire [7:0] RD_xram_69;
wire [15:0] RD_xram_69_ADDR;
wire [15:0] RD_xram_6_ADDR;
wire [7:0] RD_xram_7;
wire [7:0] RD_xram_70;
wire [15:0] RD_xram_70_ADDR;
wire [7:0] RD_xram_71;
wire [15:0] RD_xram_71_ADDR;
wire [7:0] RD_xram_72;
wire [15:0] RD_xram_72_ADDR;
wire [7:0] RD_xram_73;
wire [15:0] RD_xram_73_ADDR;
wire [7:0] RD_xram_74;
wire [15:0] RD_xram_74_ADDR;
wire [7:0] RD_xram_75;
wire [15:0] RD_xram_75_ADDR;
wire [7:0] RD_xram_76;
wire [15:0] RD_xram_76_ADDR;
wire [7:0] RD_xram_77;
wire [15:0] RD_xram_77_ADDR;
wire [7:0] RD_xram_78;
wire [15:0] RD_xram_78_ADDR;
wire [7:0] RD_xram_79;
wire [15:0] RD_xram_79_ADDR;
wire [15:0] RD_xram_7_ADDR;
wire [7:0] RD_xram_8;
wire [7:0] RD_xram_80;
wire [15:0] RD_xram_80_ADDR;
wire [15:0] RD_xram_8_ADDR;
wire [7:0] RD_xram_9;
wire [15:0] RD_xram_9_ADDR;
wire [15:0] WR_XRAM_ADDR_00;
wire [15:0] WR_XRAM_ADDR_01;
wire [15:0] WR_XRAM_ADDR_02;
wire [15:0] WR_XRAM_ADDR_03;
wire [15:0] WR_XRAM_ADDR_04;
wire [15:0] WR_XRAM_ADDR_05;
wire [15:0] WR_XRAM_ADDR_06;
wire [15:0] WR_XRAM_ADDR_07;
wire [15:0] WR_XRAM_ADDR_08;
wire [15:0] WR_XRAM_ADDR_09;
wire [15:0] WR_XRAM_ADDR_0a;
wire [15:0] WR_XRAM_ADDR_0b;
wire [15:0] WR_XRAM_ADDR_0c;
wire [15:0] WR_XRAM_ADDR_0d;
wire [15:0] WR_XRAM_ADDR_0e;
wire [15:0] WR_XRAM_ADDR_0f;
wire [15:0] WR_XRAM_ADDR_next;
wire WR_XRAM_EN_00;
wire WR_XRAM_EN_01;
wire WR_XRAM_EN_02;
wire WR_XRAM_EN_03;
wire WR_XRAM_EN_04;
wire WR_XRAM_EN_05;
wire WR_XRAM_EN_06;
wire WR_XRAM_EN_07;
wire WR_XRAM_EN_08;
wire WR_XRAM_EN_09;
wire WR_XRAM_EN_0a;
wire WR_XRAM_EN_0b;
wire WR_XRAM_EN_0c;
wire WR_XRAM_EN_0d;
wire WR_XRAM_EN_0e;
wire WR_XRAM_EN_0f;
wire WR_XRAM_EN_next;
wire [15:0] aes_addr_00;
wire [15:0] aes_addr_04;
wire [15:0] aes_addr_08;
wire [15:0] aes_addr_0c;
wire [15:0] aes_addr_next;
wire [15:0] aes_bytes_processed_00;
wire [15:0] aes_bytes_processed_01;
wire [15:0] aes_bytes_processed_02;
wire [15:0] aes_bytes_processed_03;
wire [15:0] aes_bytes_processed_04;
wire [15:0] aes_bytes_processed_05;
wire [15:0] aes_bytes_processed_06;
wire [15:0] aes_bytes_processed_07;
wire [15:0] aes_bytes_processed_08;
wire [15:0] aes_bytes_processed_09;
wire [15:0] aes_bytes_processed_0a;
wire [15:0] aes_bytes_processed_0b;
wire [15:0] aes_bytes_processed_0c;
wire [15:0] aes_bytes_processed_0d;
wire [15:0] aes_bytes_processed_0e;
wire [15:0] aes_bytes_processed_0f;
wire [15:0] aes_bytes_processed_next;
wire [127:0] aes_ctr_00;
wire [127:0] aes_ctr_04;
wire [127:0] aes_ctr_08;
wire [127:0] aes_ctr_0c;
wire [127:0] aes_ctr_next;
wire [127:0] aes_enc_data_02;
wire [127:0] aes_enc_data_06;
wire [127:0] aes_enc_data_0a;
wire [127:0] aes_enc_data_0e;
wire [127:0] aes_enc_data_next;
wire [127:0] aes_key0_00;
wire [127:0] aes_key0_04;
wire [127:0] aes_key0_08;
wire [127:0] aes_key0_0c;
wire [127:0] aes_key0_next;
wire [127:0] aes_key1_00;
wire [127:0] aes_key1_04;
wire [127:0] aes_key1_08;
wire [127:0] aes_key1_0c;
wire [127:0] aes_key1_next;
wire [15:0] aes_len_00;
wire [15:0] aes_len_04;
wire [15:0] aes_len_08;
wire [15:0] aes_len_0c;
wire [15:0] aes_len_next;
wire [127:0] aes_read_data_01;
wire [127:0] aes_read_data_05;
wire [127:0] aes_read_data_09;
wire [127:0] aes_read_data_0d;
wire [127:0] aes_read_data_next;
wire [7:0] aes_state_00;
wire [7:0] aes_state_01;
wire [7:0] aes_state_02;
wire [7:0] aes_state_03;
wire [7:0] aes_state_04;
wire [7:0] aes_state_05;
wire [7:0] aes_state_06;
wire [7:0] aes_state_07;
wire [7:0] aes_state_08;
wire [7:0] aes_state_09;
wire [7:0] aes_state_0a;
wire [7:0] aes_state_0b;
wire [7:0] aes_state_0c;
wire [7:0] aes_state_0d;
wire [7:0] aes_state_0e;
wire [7:0] aes_state_0f;
wire [7:0] aes_state_next;
wire [7:0] dataout_00;
wire [7:0] dataout_01;
wire [7:0] dataout_02;
wire [7:0] dataout_03;
wire [7:0] dataout_04;
wire [7:0] dataout_05;
wire [7:0] dataout_06;
wire [7:0] dataout_07;
wire [7:0] dataout_08;
wire [7:0] dataout_09;
wire [7:0] dataout_0a;
wire [7:0] dataout_0b;
wire [7:0] dataout_0c;
wire [7:0] dataout_0d;
wire [7:0] dataout_0e;
wire [7:0] dataout_0f;
wire [7:0] dataout_next;
wire [1:0] n0001;
wire [1:0] n0002;
wire [3:0] n0003;
wire [15:0] n0004;
wire n0005;
wire [15:0] n0006;
wire n0007;
wire [15:0] n0008;
wire n0009;
wire [15:0] n0010;
wire n0011;
wire [15:0] n0012;
wire n0013;
wire [15:0] n0014;
wire n0015;
wire [15:0] n0016;
wire n0017;
wire [15:0] n0018;
wire n0019;
wire [15:0] n0020;
wire n0021;
wire [15:0] n0022;
wire n0023;
wire [15:0] n0024;
wire n0025;
wire [15:0] n0026;
wire n0027;
wire [15:0] n0028;
wire n0029;
wire [15:0] n0030;
wire n0031;
wire [15:0] n0032;
wire [15:0] n0033;
wire [15:0] n0034;
wire [15:0] n0035;
wire n0036;
wire [15:0] n0037;
wire [15:0] n0038;
wire [15:0] n0039;
wire [15:0] n0040;
wire [15:0] n0041;
wire [15:0] n0042;
wire [15:0] n0043;
wire [15:0] n0044;
wire [15:0] n0045;
wire [15:0] n0046;
wire [15:0] n0047;
wire [15:0] n0048;
wire [15:0] n0049;
wire [15:0] n0050;
wire [15:0] n0051;
wire [15:0] n0052;
wire [15:0] n0053;
wire [15:0] n0054;
wire [15:0] n0055;
wire [15:0] n0056;
wire [15:0] n0057;
wire [15:0] n0058;
wire [15:0] n0059;
wire [15:0] n0060;
wire [15:0] n0061;
wire [15:0] n0062;
wire [15:0] n0063;
wire [15:0] n0064;
wire [15:0] n0065;
wire [15:0] n0066;
wire [15:0] n0067;
wire [15:0] n0068;
wire [15:0] n0069;
wire [15:0] n0070;
wire [15:0] n0071;
wire [15:0] n0072;
wire [15:0] n0073;
wire [15:0] n0074;
wire [15:0] n0075;
wire [15:0] n0076;
wire [15:0] n0077;
wire [15:0] n0078;
wire [15:0] n0079;
wire [15:0] n0080;
wire [15:0] n0081;
wire [15:0] n0082;
wire [15:0] n0083;
wire [15:0] n0084;
wire [15:0] n0085;
wire [15:0] n0086;
wire [15:0] n0087;
wire [15:0] n0088;
wire [15:0] n0089;
wire [15:0] n0090;
wire [15:0] n0091;
wire [15:0] n0092;
wire [15:0] n0093;
wire [15:0] n0094;
wire [15:0] n0095;
wire [15:0] n0096;
wire [15:0] n0097;
wire [15:0] n0098;
wire [15:0] n0099;
wire [15:0] n0100;
wire [15:0] n0101;
wire [15:0] n0102;
wire [15:0] n0103;
wire [15:0] n0104;
wire [15:0] n0105;
wire [15:0] n0106;
wire [15:0] n0107;
wire [15:0] n0108;
wire [15:0] n0109;
wire [15:0] n0110;
wire [15:0] n0111;
wire [15:0] n0112;
wire [15:0] n0113;
wire [15:0] n0114;
wire [15:0] n0115;
wire [15:0] n0116;
wire [15:0] n0117;
wire [15:0] n0118;
wire [15:0] n0119;
wire [15:0] n0120;
wire [15:0] n0121;
wire [15:0] n0122;
wire [15:0] n0123;
wire [15:0] n0124;
wire [15:0] n0125;
wire [15:0] n0126;
wire [15:0] n0127;
wire [15:0] n0128;
wire [15:0] n0129;
wire [15:0] n0130;
wire [15:0] n0131;
wire [15:0] n0132;
wire [15:0] n0133;
wire [15:0] n0134;
wire [15:0] n0135;
wire [15:0] n0136;
wire [15:0] n0137;
wire [15:0] n0138;
wire [15:0] n0139;
wire [15:0] n0140;
wire [15:0] n0141;
wire [15:0] n0142;
wire [15:0] n0143;
wire [15:0] n0144;
wire [15:0] n0145;
wire [15:0] n0146;
wire [15:0] n0147;
wire [15:0] n0148;
wire [15:0] n0149;
wire [15:0] n0150;
wire [15:0] n0151;
wire [15:0] n0152;
wire [15:0] n0153;
wire [15:0] n0154;
wire [15:0] n0155;
wire [15:0] n0156;
wire [15:0] n0157;
wire [15:0] n0158;
wire [15:0] n0159;
wire [15:0] n0160;
wire [15:0] n0161;
wire [15:0] n0162;
wire [15:0] n0163;
wire [15:0] n0164;
wire [15:0] n0165;
wire [15:0] n0166;
wire [15:0] n0167;
wire [15:0] n0168;
wire [15:0] n0169;
wire [15:0] n0170;
wire [15:0] n0171;
wire [15:0] n0172;
wire [15:0] n0173;
wire [15:0] n0174;
wire [15:0] n0175;
wire [15:0] n0176;
wire [15:0] n0177;
wire [15:0] n0178;
wire [15:0] n0179;
wire [15:0] n0180;
wire [15:0] n0181;
wire [15:0] n0182;
wire [15:0] n0183;
wire [15:0] n0184;
wire [15:0] n0185;
wire [15:0] n0186;
wire [15:0] n0187;
wire [15:0] n0188;
wire [15:0] n0189;
wire [15:0] n0190;
wire [15:0] n0191;
wire [15:0] n0192;
wire [15:0] n0193;
wire [15:0] n0194;
wire [15:0] n0195;
wire [15:0] n0196;
wire [15:0] n0197;
wire [15:0] n0198;
wire [15:0] n0199;
wire [15:0] n0200;
wire [15:0] n0201;
wire [15:0] n0202;
wire [15:0] n0203;
wire [15:0] n0204;
wire [15:0] n0205;
wire [15:0] n0206;
wire [15:0] n0207;
wire [15:0] n0208;
wire [15:0] n0209;
wire [15:0] n0210;
wire [15:0] n0211;
wire [15:0] n0212;
wire [15:0] n0213;
wire [15:0] n0214;
wire [15:0] n0215;
wire [15:0] n0216;
wire [15:0] n0217;
wire [15:0] n0218;
wire [15:0] n0219;
wire [15:0] n0220;
wire [15:0] n0221;
wire [15:0] n0222;
wire [15:0] n0223;
wire [15:0] n0224;
wire [15:0] n0225;
wire [15:0] n0226;
wire [15:0] n0227;
wire [15:0] n0228;
wire [15:0] n0229;
wire [15:0] n0230;
wire [15:0] n0231;
wire [15:0] n0232;
wire [15:0] n0233;
wire [15:0] n0234;
wire [15:0] n0235;
wire [15:0] n0236;
wire [15:0] n0237;
wire [15:0] n0238;
wire [15:0] n0239;
wire [15:0] n0240;
wire [15:0] n0241;
wire [15:0] n0242;
wire [15:0] n0243;
wire [15:0] n0244;
wire [15:0] n0245;
wire [15:0] n0246;
wire [15:0] n0247;
wire [15:0] n0248;
wire [15:0] n0249;
wire [15:0] n0250;
wire [15:0] n0251;
wire [15:0] n0252;
wire [15:0] n0253;
wire [15:0] n0254;
wire [15:0] n0255;
wire [15:0] n0256;
wire [15:0] n0257;
wire [15:0] n0258;
wire [15:0] n0259;
wire [15:0] n0260;
wire [15:0] n0261;
wire [15:0] n0262;
wire [15:0] n0263;
wire [15:0] n0264;
wire [15:0] n0265;
wire [15:0] n0266;
wire [15:0] n0267;
wire [15:0] n0268;
wire [15:0] n0269;
wire [15:0] n0270;
wire [15:0] n0271;
wire [15:0] n0272;
wire [15:0] n0273;
wire [15:0] n0274;
wire [15:0] n0275;
wire [15:0] n0276;
wire [15:0] n0277;
wire [15:0] n0278;
wire [15:0] n0279;
wire [15:0] n0280;
wire [15:0] n0281;
wire [15:0] n0282;
wire [15:0] n0283;
wire [15:0] n0284;
wire [15:0] n0285;
wire [15:0] n0286;
wire [15:0] n0287;
wire [15:0] n0288;
wire [15:0] n0289;
wire [15:0] n0290;
wire [15:0] n0291;
wire [15:0] n0292;
wire [15:0] n0293;
wire [15:0] n0294;
wire [15:0] n0295;
wire [15:0] n0296;
wire [15:0] n0297;
wire [15:0] n0298;
wire [15:0] n0299;
wire [15:0] n0300;
wire [15:0] n0301;
wire [15:0] n0302;
wire [15:0] n0303;
wire [15:0] n0304;
wire [15:0] n0305;
wire [15:0] n0306;
wire [15:0] n0307;
wire [15:0] n0308;
wire [15:0] n0309;
wire [15:0] n0310;
wire [15:0] n0311;
wire [15:0] n0312;
wire [15:0] n0313;
wire [15:0] n0314;
wire [15:0] n0315;
wire [15:0] n0316;
wire [15:0] n0317;
wire [15:0] n0318;
wire [15:0] n0319;
wire [15:0] n0320;
wire [15:0] n0321;
wire [15:0] n0322;
wire [15:0] n0323;
wire [15:0] n0324;
wire [15:0] n0325;
wire [15:0] n0326;
wire [15:0] n0327;
wire [15:0] n0328;
wire [15:0] n0329;
wire [15:0] n0330;
wire [15:0] n0331;
wire [15:0] n0332;
wire [15:0] n0333;
wire [15:0] n0334;
wire [15:0] n0335;
wire [15:0] n0336;
wire [15:0] n0337;
wire [15:0] n0338;
wire [15:0] n0339;
wire [15:0] n0340;
wire [15:0] n0341;
wire [15:0] n0342;
wire [15:0] n0343;
wire [15:0] n0344;
wire [15:0] n0345;
wire [15:0] n0346;
wire [15:0] n0347;
wire [15:0] n0348;
wire [15:0] n0349;
wire [15:0] n0350;
wire [15:0] n0351;
wire [15:0] n0352;
wire [15:0] n0353;
wire [15:0] n0354;
wire [15:0] n0355;
wire [15:0] n0356;
wire [15:0] n0357;
wire [15:0] n0358;
wire [15:0] n0359;
wire [15:0] n0360;
wire [15:0] n0361;
wire [15:0] n0362;
wire [15:0] n0363;
wire [15:0] n0364;
wire [15:0] n0365;
wire [15:0] n0366;
wire [15:0] n0367;
wire [15:0] n0368;
wire [15:0] n0369;
wire [15:0] n0370;
wire [15:0] n0371;
wire [15:0] n0372;
wire [15:0] n0373;
wire [15:0] n0374;
wire [15:0] n0375;
wire [15:0] n0376;
wire [15:0] n0377;
wire [15:0] n0378;
wire [15:0] n0379;
wire [15:0] n0380;
wire [15:0] n0381;
wire [15:0] n0382;
wire [15:0] n0383;
wire [15:0] n0384;
wire [15:0] n0385;
wire [15:0] n0386;
wire [15:0] n0387;
wire [15:0] n0388;
wire [15:0] n0389;
wire [15:0] n0390;
wire [15:0] n0391;
wire [15:0] n0392;
wire [15:0] n0393;
wire [15:0] n0394;
wire [15:0] n0395;
wire [15:0] n0396;
wire [15:0] n0397;
wire [15:0] n0398;
wire [15:0] n0399;
wire [15:0] n0400;
wire [15:0] n0401;
wire [15:0] n0402;
wire [15:0] n0403;
wire [15:0] n0404;
wire [15:0] n0405;
wire [15:0] n0406;
wire [15:0] n0407;
wire [15:0] n0408;
wire [15:0] n0409;
wire [15:0] n0410;
wire [15:0] n0411;
wire [15:0] n0412;
wire [15:0] n0413;
wire [15:0] n0414;
wire [15:0] n0415;
wire [15:0] n0416;
wire [15:0] n0417;
wire [15:0] n0418;
wire [15:0] n0419;
wire [15:0] n0420;
wire [15:0] n0421;
wire [15:0] n0422;
wire [15:0] n0423;
wire [15:0] n0424;
wire [15:0] n0425;
wire [15:0] n0426;
wire [15:0] n0427;
wire [15:0] n0428;
wire [15:0] n0429;
wire [15:0] n0430;
wire [15:0] n0431;
wire [15:0] n0432;
wire [15:0] n0433;
wire [15:0] n0434;
wire [15:0] n0435;
wire [15:0] n0436;
wire [15:0] n0437;
wire [15:0] n0438;
wire [15:0] n0439;
wire [15:0] n0440;
wire [15:0] n0441;
wire [15:0] n0442;
wire [15:0] n0443;
wire [15:0] n0444;
wire [15:0] n0445;
wire [15:0] n0446;
wire [15:0] n0447;
wire [15:0] n0448;
wire [15:0] n0449;
wire [15:0] n0450;
wire [15:0] n0451;
wire [15:0] n0452;
wire [15:0] n0453;
wire [15:0] n0454;
wire [15:0] n0455;
wire [15:0] n0456;
wire [15:0] n0457;
wire [15:0] n0458;
wire [15:0] n0459;
wire [15:0] n0460;
wire [15:0] n0461;
wire [15:0] n0462;
wire [15:0] n0463;
wire [15:0] n0464;
wire [15:0] n0465;
wire [15:0] n0466;
wire [15:0] n0467;
wire [15:0] n0468;
wire [15:0] n0469;
wire [15:0] n0470;
wire [15:0] n0471;
wire [15:0] n0472;
wire [15:0] n0473;
wire [15:0] n0474;
wire [15:0] n0475;
wire [15:0] n0476;
wire [15:0] n0477;
wire [15:0] n0478;
wire [15:0] n0479;
wire [15:0] n0480;
wire [15:0] n0481;
wire [15:0] n0482;
wire [15:0] n0483;
wire [15:0] n0484;
wire [15:0] n0485;
wire [15:0] n0486;
wire [15:0] n0487;
wire [15:0] n0488;
wire [15:0] n0489;
wire [15:0] n0490;
wire [15:0] n0491;
wire [15:0] n0492;
wire [15:0] n0493;
wire [15:0] n0494;
wire [15:0] n0495;
wire [15:0] n0496;
wire [15:0] n0497;
wire [15:0] n0498;
wire n0499;
wire [15:0] n0500;
wire n0501;
wire n0502;
wire [15:0] n0503;
wire n0504;
wire [1:0] n0505;
wire [1:0] n0506;
wire n0507;
wire n0508;
wire [15:0] n0509;
wire [14:0] n0510;
wire [0:0] n0511;
wire [15:0] n0512;
wire n0513;
wire n0514;
wire [0:0] n0515;
wire n0516;
wire [7:0] n0517;
wire [7:0] n0518;
wire [7:0] n0519;
wire [15:0] n0520;
wire n0521;
wire n0522;
wire [7:0] n0523;
wire [7:0] n0524;
wire [7:0] n0525;
wire [15:0] n0526;
wire [11:0] n0527;
wire [3:0] n0528;
wire [15:0] n0529;
wire n0530;
wire n0531;
wire [3:0] n0532;
wire n0533;
wire [7:0] n0534;
wire [3:0] n0535;
wire n0536;
wire [7:0] n0537;
wire [3:0] n0538;
wire n0539;
wire [7:0] n0540;
wire [3:0] n0541;
wire n0542;
wire [7:0] n0543;
wire [3:0] n0544;
wire n0545;
wire [7:0] n0546;
wire [3:0] n0547;
wire n0548;
wire [7:0] n0549;
wire [3:0] n0550;
wire n0551;
wire [7:0] n0552;
wire [3:0] n0553;
wire n0554;
wire [7:0] n0555;
wire [3:0] n0556;
wire n0557;
wire [7:0] n0558;
wire [3:0] n0559;
wire n0560;
wire [7:0] n0561;
wire [3:0] n0562;
wire n0563;
wire [7:0] n0564;
wire [3:0] n0565;
wire n0566;
wire [7:0] n0567;
wire [3:0] n0568;
wire n0569;
wire [7:0] n0570;
wire [3:0] n0571;
wire n0572;
wire [7:0] n0573;
wire [3:0] n0574;
wire n0575;
wire [7:0] n0576;
wire [7:0] n0577;
wire [7:0] n0578;
wire [7:0] n0579;
wire [7:0] n0580;
wire [7:0] n0581;
wire [7:0] n0582;
wire [7:0] n0583;
wire [7:0] n0584;
wire [7:0] n0585;
wire [7:0] n0586;
wire [7:0] n0587;
wire [7:0] n0588;
wire [7:0] n0589;
wire [7:0] n0590;
wire [7:0] n0591;
wire [7:0] n0592;
wire [15:0] n0593;
wire n0594;
wire n0595;
wire [7:0] n0596;
wire [7:0] n0597;
wire [7:0] n0598;
wire [7:0] n0599;
wire [7:0] n0600;
wire [7:0] n0601;
wire [7:0] n0602;
wire [7:0] n0603;
wire [7:0] n0604;
wire [7:0] n0605;
wire [7:0] n0606;
wire [7:0] n0607;
wire [7:0] n0608;
wire [7:0] n0609;
wire [7:0] n0610;
wire [7:0] n0611;
wire [7:0] n0612;
wire [7:0] n0613;
wire [7:0] n0614;
wire [7:0] n0615;
wire [7:0] n0616;
wire [7:0] n0617;
wire [7:0] n0618;
wire [7:0] n0619;
wire [7:0] n0620;
wire [7:0] n0621;
wire [7:0] n0622;
wire [7:0] n0623;
wire [7:0] n0624;
wire [7:0] n0625;
wire [7:0] n0626;
wire [15:0] n0627;
wire n0628;
wire n0629;
wire [7:0] n0630;
wire [7:0] n0631;
wire [7:0] n0632;
wire [7:0] n0633;
wire [7:0] n0634;
wire [7:0] n0635;
wire [7:0] n0636;
wire [7:0] n0637;
wire [7:0] n0638;
wire [7:0] n0639;
wire [7:0] n0640;
wire [7:0] n0641;
wire [7:0] n0642;
wire [7:0] n0643;
wire [7:0] n0644;
wire [7:0] n0645;
wire [7:0] n0646;
wire [7:0] n0647;
wire [7:0] n0648;
wire [7:0] n0649;
wire [7:0] n0650;
wire [7:0] n0651;
wire [7:0] n0652;
wire [7:0] n0653;
wire [7:0] n0654;
wire [7:0] n0655;
wire [7:0] n0656;
wire [7:0] n0657;
wire [7:0] n0658;
wire [7:0] n0659;
wire [7:0] n0660;
wire [7:0] n0661;
wire [7:0] n0662;
wire [7:0] n0663;
wire [7:0] n0664;
wire [7:0] n0665;
wire [7:0] n0666;
wire [7:0] n0667;
wire [15:0] n0668;
wire n0669;
wire [15:0] n0670;
wire n0671;
wire n0672;
wire n0673;
wire n0674;
wire [15:0] n0675;
wire n0676;
wire n0677;
wire [7:0] n0678;
wire [7:0] n0679;
wire [7:0] n0680;
wire [15:0] n0681;
wire n0682;
wire n0683;
wire [7:0] n0684;
wire [7:0] n0685;
wire [7:0] n0686;
wire [15:0] n0687;
wire n0688;
wire n0689;
wire [7:0] n0690;
wire [7:0] n0691;
wire [7:0] n0692;
wire [7:0] n0693;
wire [7:0] n0694;
wire [7:0] n0695;
wire [7:0] n0696;
wire [7:0] n0697;
wire [7:0] n0698;
wire [7:0] n0699;
wire [1:0] n0700;
wire n0701;
wire n0702;
wire [15:0] n0703;
wire [15:0] n0704;
wire [15:0] n0705;
wire [15:0] n0706;
wire n0707;
wire n0708;
wire n0709;
wire [15:0] n0710;
wire [15:0] n0711;
wire [15:0] n0712;
wire [15:0] n0713;
wire n0714;
wire [119:0] n0715;
wire [127:0] n0716;
wire [111:0] n0717;
wire [127:0] n0718;
wire [103:0] n0719;
wire [15:0] n0720;
wire [127:0] n0721;
wire [95:0] n0722;
wire [23:0] n0723;
wire [127:0] n0724;
wire [87:0] n0725;
wire [31:0] n0726;
wire [127:0] n0727;
wire [79:0] n0728;
wire [39:0] n0729;
wire [127:0] n0730;
wire [71:0] n0731;
wire [47:0] n0732;
wire [127:0] n0733;
wire [63:0] n0734;
wire [55:0] n0735;
wire [127:0] n0736;
wire [55:0] n0737;
wire [63:0] n0738;
wire [127:0] n0739;
wire [47:0] n0740;
wire [71:0] n0741;
wire [127:0] n0742;
wire [39:0] n0743;
wire [79:0] n0744;
wire [127:0] n0745;
wire [31:0] n0746;
wire [87:0] n0747;
wire [127:0] n0748;
wire [23:0] n0749;
wire [95:0] n0750;
wire [127:0] n0751;
wire [15:0] n0752;
wire [103:0] n0753;
wire [127:0] n0754;
wire [111:0] n0755;
wire [127:0] n0756;
wire [119:0] n0757;
wire [127:0] n0758;
wire [127:0] n0759;
wire [127:0] n0760;
wire [127:0] n0761;
wire [127:0] n0762;
wire [127:0] n0763;
wire [127:0] n0764;
wire [127:0] n0765;
wire [127:0] n0766;
wire [127:0] n0767;
wire [127:0] n0768;
wire [127:0] n0769;
wire [127:0] n0770;
wire [127:0] n0771;
wire [127:0] n0772;
wire [127:0] n0773;
wire [127:0] n0774;
wire [0:0] n0775;
wire [0:0] n0776;
wire n0777;
wire n0778;
wire n0779;
wire [15:0] n0780;
wire n0781;
wire [15:0] n0782;
wire [15:0] n0783;
wire [15:0] n0784;
wire [15:0] n0785;
wire n0786;
wire [119:0] n0787;
wire [127:0] n0788;
wire [111:0] n0789;
wire [127:0] n0790;
wire [103:0] n0791;
wire [15:0] n0792;
wire [127:0] n0793;
wire [95:0] n0794;
wire [23:0] n0795;
wire [127:0] n0796;
wire [87:0] n0797;
wire [31:0] n0798;
wire [127:0] n0799;
wire [79:0] n0800;
wire [39:0] n0801;
wire [127:0] n0802;
wire [71:0] n0803;
wire [47:0] n0804;
wire [127:0] n0805;
wire [63:0] n0806;
wire [55:0] n0807;
wire [127:0] n0808;
wire [55:0] n0809;
wire [63:0] n0810;
wire [127:0] n0811;
wire [47:0] n0812;
wire [71:0] n0813;
wire [127:0] n0814;
wire [39:0] n0815;
wire [79:0] n0816;
wire [127:0] n0817;
wire [31:0] n0818;
wire [87:0] n0819;
wire [127:0] n0820;
wire [23:0] n0821;
wire [95:0] n0822;
wire [127:0] n0823;
wire [15:0] n0824;
wire [103:0] n0825;
wire [127:0] n0826;
wire [111:0] n0827;
wire [127:0] n0828;
wire [119:0] n0829;
wire [127:0] n0830;
wire [127:0] n0831;
wire [127:0] n0832;
wire [127:0] n0833;
wire [127:0] n0834;
wire [127:0] n0835;
wire [127:0] n0836;
wire [127:0] n0837;
wire [127:0] n0838;
wire [127:0] n0839;
wire [127:0] n0840;
wire [127:0] n0841;
wire [127:0] n0842;
wire [127:0] n0843;
wire [127:0] n0844;
wire [127:0] n0845;
wire [127:0] n0846;
wire n0847;
wire [119:0] n0848;
wire [127:0] n0849;
wire [111:0] n0850;
wire [127:0] n0851;
wire [103:0] n0852;
wire [15:0] n0853;
wire [127:0] n0854;
wire [95:0] n0855;
wire [23:0] n0856;
wire [127:0] n0857;
wire [87:0] n0858;
wire [31:0] n0859;
wire [127:0] n0860;
wire [79:0] n0861;
wire [39:0] n0862;
wire [127:0] n0863;
wire [71:0] n0864;
wire [47:0] n0865;
wire [127:0] n0866;
wire [63:0] n0867;
wire [55:0] n0868;
wire [127:0] n0869;
wire [55:0] n0870;
wire [63:0] n0871;
wire [127:0] n0872;
wire [47:0] n0873;
wire [71:0] n0874;
wire [127:0] n0875;
wire [39:0] n0876;
wire [79:0] n0877;
wire [127:0] n0878;
wire [31:0] n0879;
wire [87:0] n0880;
wire [127:0] n0881;
wire [23:0] n0882;
wire [95:0] n0883;
wire [127:0] n0884;
wire [15:0] n0885;
wire [103:0] n0886;
wire [127:0] n0887;
wire [111:0] n0888;
wire [127:0] n0889;
wire [119:0] n0890;
wire [127:0] n0891;
wire [127:0] n0892;
wire [127:0] n0893;
wire [127:0] n0894;
wire [127:0] n0895;
wire [127:0] n0896;
wire [127:0] n0897;
wire [127:0] n0898;
wire [127:0] n0899;
wire [127:0] n0900;
wire [127:0] n0901;
wire [127:0] n0902;
wire [127:0] n0903;
wire [127:0] n0904;
wire [127:0] n0905;
wire [127:0] n0906;
wire [127:0] n0907;
wire n0908;
wire [15:0] n0909;
wire [15:0] n0910;
wire [15:0] n0911;
wire [15:0] n0912;
wire n0913;
wire n0914;
wire n0915;
wire [7:0] n0916;
wire [7:0] n0917;
wire [15:0] n0918;
wire n0919;
wire [15:0] n0920;
wire [15:0] n0921;
wire [15:0] n0922;
wire [15:0] n0923;
wire n0924;
wire [159:0] n0925;
wire [159:0] n0926;
wire [7:0] n0927;
wire n0928;
wire [0:0] n0929;
wire n0930;
wire [159:0] n0931;
wire [159:0] n0932;
wire [159:0] n0933;
wire [159:0] n0934;
wire [7:0] n0935;
wire n0936;
wire n0937;
wire n0938;
wire n0939;
wire [15:0] n0940;
wire n0941;
wire n0942;
wire [7:0] n0943;
wire [15:0] n0944;
wire n0945;
wire n0946;
wire [7:0] n0947;
wire [7:0] n0948;
wire [7:0] n0949;
wire [15:0] n0950;
wire n0951;
wire n0952;
wire [15:0] n0953;
wire [0:0] n0954;
wire n0955;
wire [127:0] n0956;
wire [127:0] n0957;
wire [159:0] n0958;
wire [159:0] n0959;
wire [159:0] n0960;
wire [159:0] n0961;
wire [7:0] n0962;
wire [7:0] n0963;
wire [7:0] n0964;
wire [7:0] n0965;
wire [127:0] n0966;
wire [127:0] n0967;
wire [159:0] n0968;
wire [159:0] n0969;
wire [159:0] n0970;
wire [159:0] n0971;
wire [15:0] n0972;
wire [15:0] n0973;
wire [15:0] n0974;
wire n0975;
wire n0976;
wire [7:0] n0977;
wire [7:0] n0978;
wire [7:0] n0979;
wire n0980;
wire [7:0] n0981;
wire [7:0] n0982;
wire [159:0] n0983;
wire [159:0] n0984;
wire [159:0] n0985;
wire [159:0] n0986;
wire n0987;
wire n0988;
wire n0989;
wire n0990;
wire n0991;
wire n0992;
wire n0993;
wire n0994;
wire n0995;
wire n0996;
wire n0997;
wire n0998;
wire n0999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire [15:0] n1102;
wire [15:0] n1103;
wire [15:0] n1104;
wire [15:0] n1105;
wire [15:0] n1106;
wire [15:0] n1107;
wire [15:0] n1108;
wire [15:0] n1109;
wire [15:0] n1110;
wire [15:0] n1111;
wire [15:0] n1112;
wire [15:0] n1113;
wire [15:0] n1114;
wire [15:0] n1115;
wire [15:0] n1116;
wire [15:0] n1117;
wire [15:0] n1118;
wire [15:0] n1119;
wire [15:0] n1120;
wire [15:0] n1121;
wire [15:0] n1122;
wire [15:0] n1123;
wire [15:0] n1124;
wire [15:0] n1125;
wire [15:0] n1126;
wire [15:0] n1127;
wire [15:0] n1128;
wire [15:0] n1129;
wire [15:0] n1130;
wire [15:0] n1131;
wire [15:0] n1132;
wire [15:0] n1133;
wire [15:0] n1134;
wire [15:0] n1135;
wire [15:0] n1136;
wire [15:0] n1137;
wire [15:0] n1138;
wire [15:0] n1139;
wire [15:0] n1140;
wire [15:0] n1141;
wire [15:0] n1142;
wire [15:0] n1143;
wire [15:0] n1144;
wire [15:0] n1145;
wire [15:0] n1146;
wire [15:0] n1147;
wire [15:0] n1148;
wire [15:0] n1149;
wire [15:0] n1150;
wire [15:0] n1151;
wire [15:0] n1152;
wire [15:0] n1153;
wire [15:0] n1154;
wire [15:0] n1155;
wire [15:0] n1156;
wire [15:0] n1157;
wire [15:0] n1158;
wire [15:0] n1159;
wire [15:0] n1160;
wire [15:0] n1161;
wire [15:0] n1162;
wire [15:0] n1163;
wire [15:0] n1164;
wire [15:0] n1165;
wire [15:0] n1166;
wire [15:0] n1167;
wire [15:0] n1168;
wire [15:0] n1169;
wire [15:0] n1170;
wire [15:0] n1171;
wire [15:0] n1172;
wire [15:0] n1173;
wire [15:0] n1174;
wire [15:0] n1175;
wire [15:0] n1176;
wire [15:0] n1177;
wire [15:0] n1178;
wire [15:0] n1179;
wire [15:0] n1180;
wire [15:0] n1181;
wire [15:0] n1182;
wire [15:0] n1183;
wire [15:0] n1184;
wire [15:0] n1185;
wire [15:0] n1186;
wire [15:0] n1187;
wire [15:0] n1188;
wire [15:0] n1189;
wire [15:0] n1190;
wire [15:0] n1191;
wire [15:0] n1192;
wire [15:0] n1193;
wire [15:0] n1194;
wire [15:0] n1195;
wire [15:0] n1196;
wire [15:0] n1197;
wire [15:0] n1198;
wire [15:0] n1199;
wire [15:0] n1200;
wire [15:0] n1201;
wire [15:0] n1202;
wire [15:0] n1203;
wire [15:0] n1204;
wire [15:0] n1205;
wire [15:0] n1206;
wire [15:0] n1207;
wire [15:0] n1208;
wire [15:0] n1209;
wire [15:0] n1210;
wire [15:0] n1211;
wire [15:0] n1212;
wire [15:0] n1213;
wire [15:0] n1214;
wire [15:0] n1215;
wire [15:0] n1216;
wire [15:0] n1217;
wire [15:0] n1218;
wire [15:0] n1219;
wire [15:0] n1220;
wire [15:0] n1221;
wire [15:0] n1222;
wire [15:0] n1223;
wire [15:0] n1224;
wire [15:0] n1225;
wire [15:0] n1226;
wire n1227;
wire n1228;
wire [7:0] n1229;
wire [15:0] n1230;
wire n1231;
wire n1232;
wire [7:0] n1233;
wire [7:0] n1234;
wire [7:0] n1235;
wire [159:0] n1236;
wire [159:0] n1237;
wire [159:0] n1238;
wire [159:0] n1239;
wire [511:0] n1240;
wire [511:0] n1241;
wire [7:0] n1242;
wire [7:0] n1243;
wire [159:0] n1244;
wire [159:0] n1245;
wire [159:0] n1246;
wire [159:0] n1247;
wire [511:0] n1248;
wire [511:0] n1249;
wire [159:0] n1250;
wire [159:0] n1251;
wire [159:0] n1252;
wire [159:0] n1253;
wire [127:0] n1254;
wire [127:0] n1255;
wire [159:0] n1256;
wire [159:0] n1257;
wire [159:0] n1258;
wire [159:0] n1259;
wire [7:0] n1260;
wire [15:0] n1261;
wire [15:0] n1262;
wire [15:0] n1263;
wire n1264;
wire [7:0] n1265;
wire [7:0] n1266;
wire [159:0] n1267;
wire [159:0] n1268;
wire [159:0] n1269;
wire [159:0] n1270;
wire [159:0] n1271;
wire [159:0] n1272;
wire [159:0] n1273;
wire [159:0] n1274;
wire [159:0] n1275;
wire [159:0] n1276;
wire [159:0] n1277;
wire [159:0] n1278;
wire [127:0] n1279;
wire [127:0] n1280;
wire [159:0] n1281;
wire [159:0] n1282;
wire [159:0] n1283;
wire [159:0] n1284;
wire [159:0] n1285;
wire [159:0] n1286;
wire [159:0] n1287;
wire [159:0] n1288;
wire [7:0] n1289;
wire [127:0] n1290;
wire [127:0] n1291;
wire [7:0] n1292;
wire [7:0] n1293;
wire [7:0] n1294;
wire [159:0] n1295;
wire [159:0] n1296;
wire [159:0] n1297;
wire [159:0] n1298;
wire [159:0] n1299;
wire [159:0] n1300;
wire [159:0] n1301;
wire [159:0] n1302;
wire [127:0] n1303;
wire [127:0] n1304;
wire [159:0] n1305;
wire [159:0] n1306;
wire [159:0] n1307;
wire [159:0] n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire [3:0] n1324;
wire n1325;
wire [15:0] sha_bytes_processed_00;
wire [15:0] sha_bytes_processed_01;
wire [15:0] sha_bytes_processed_02;
wire [15:0] sha_bytes_processed_03;
wire [15:0] sha_bytes_processed_04;
wire [15:0] sha_bytes_processed_05;
wire [15:0] sha_bytes_processed_06;
wire [15:0] sha_bytes_processed_07;
wire [15:0] sha_bytes_processed_08;
wire [15:0] sha_bytes_processed_09;
wire [15:0] sha_bytes_processed_0a;
wire [15:0] sha_bytes_processed_0b;
wire [15:0] sha_bytes_processed_0c;
wire [15:0] sha_bytes_processed_0d;
wire [15:0] sha_bytes_processed_0e;
wire [15:0] sha_bytes_processed_0f;
wire [15:0] sha_bytes_processed_next;
wire [159:0] sha_digest_00;
wire [159:0] sha_digest_01;
wire [159:0] sha_digest_02;
wire [159:0] sha_digest_03;
wire [159:0] sha_digest_04;
wire [159:0] sha_digest_05;
wire [159:0] sha_digest_06;
wire [159:0] sha_digest_07;
wire [159:0] sha_digest_08;
wire [159:0] sha_digest_09;
wire [159:0] sha_digest_0a;
wire [159:0] sha_digest_0b;
wire [159:0] sha_digest_0c;
wire [159:0] sha_digest_0d;
wire [159:0] sha_digest_0e;
wire [159:0] sha_digest_0f;
wire [159:0] sha_digest_next;
wire [15:0] sha_len_00;
wire [15:0] sha_len_01;
wire [15:0] sha_len_02;
wire [15:0] sha_len_03;
wire [15:0] sha_len_next;
wire [15:0] sha_rdaddr_00;
wire [15:0] sha_rdaddr_01;
wire [15:0] sha_rdaddr_02;
wire [15:0] sha_rdaddr_03;
wire [15:0] sha_rdaddr_next;
wire [511:0] sha_read_data_04;
wire [511:0] sha_read_data_05;
wire [511:0] sha_read_data_06;
wire [511:0] sha_read_data_07;
wire [511:0] sha_read_data_next;
wire [7:0] sha_state_00;
wire [7:0] sha_state_01;
wire [7:0] sha_state_02;
wire [7:0] sha_state_03;
wire [7:0] sha_state_04;
wire [7:0] sha_state_05;
wire [7:0] sha_state_06;
wire [7:0] sha_state_07;
wire [7:0] sha_state_08;
wire [7:0] sha_state_09;
wire [7:0] sha_state_0a;
wire [7:0] sha_state_0b;
wire [7:0] sha_state_0c;
wire [7:0] sha_state_0d;
wire [7:0] sha_state_0e;
wire [7:0] sha_state_0f;
wire [7:0] sha_state_next;
wire [15:0] sha_wraddr_00;
wire [15:0] sha_wraddr_01;
wire [15:0] sha_wraddr_02;
wire [15:0] sha_wraddr_03;
wire [15:0] sha_wraddr_next;


// port: xram->RD_xram_0
// port: xram->RD_xram_1
// port: xram->RD_xram_2
// port: xram->RD_xram_3
// port: xram->RD_xram_4
// port: xram->RD_xram_5
// port: xram->RD_xram_6
// port: xram->RD_xram_7
// port: xram->RD_xram_8
// port: xram->RD_xram_9
// port: xram->RD_xram_10
// port: xram->RD_xram_11
// port: xram->RD_xram_12
// port: xram->RD_xram_13
// port: xram->RD_xram_14
// port: xram->RD_xram_15
// port: xram->RD_xram_16
// port: xram->RD_xram_17
// port: xram->RD_xram_18
// port: xram->RD_xram_19
// port: xram->RD_xram_20
// port: xram->RD_xram_21
// port: xram->RD_xram_22
// port: xram->RD_xram_23
// port: xram->RD_xram_24
// port: xram->RD_xram_25
// port: xram->RD_xram_26
// port: xram->RD_xram_27
// port: xram->RD_xram_28
// port: xram->RD_xram_29
// port: xram->RD_xram_30
// port: xram->RD_xram_31
// port: xram->RD_xram_32
// port: xram->RD_xram_33
// port: xram->RD_xram_34
// port: xram->RD_xram_35
// port: xram->RD_xram_36
// port: xram->RD_xram_37
// port: xram->RD_xram_38
// port: xram->RD_xram_39
// port: xram->RD_xram_40
// port: xram->RD_xram_41
// port: xram->RD_xram_42
// port: xram->RD_xram_43
// port: xram->RD_xram_44
// port: xram->RD_xram_45
// port: xram->RD_xram_46
// port: xram->RD_xram_47
// port: xram->RD_xram_48
// port: xram->RD_xram_49
// port: xram->RD_xram_50
// port: xram->RD_xram_51
// port: xram->RD_xram_52
// port: xram->RD_xram_53
// port: xram->RD_xram_54
// port: xram->RD_xram_55
// port: xram->RD_xram_56
// port: xram->RD_xram_57
// port: xram->RD_xram_58
// port: xram->RD_xram_59
// port: xram->RD_xram_60
// port: xram->RD_xram_61
// port: xram->RD_xram_62
// port: xram->RD_xram_63
// port: xram->RD_xram_64
// port: xram->RD_xram_65
// port: xram->RD_xram_66
// port: xram->RD_xram_67
// port: xram->RD_xram_68
// port: xram->RD_xram_69
// port: xram->RD_xram_70
// port: xram->RD_xram_71
// port: xram->RD_xram_72
// port: xram->RD_xram_73
// port: xram->RD_xram_74
// port: xram->RD_xram_75
// port: xram->RD_xram_76
// port: xram->RD_xram_77
// port: xram->RD_xram_78
// port: xram->RD_xram_79
// port: xram->RD_xram_80
// RD_xram_0_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 0 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 2 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 3 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 8 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 10 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 11 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 12 16)) addrin (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 13 16)) (add aes_addr (add aes_bytes_processed (bv 15 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 14 16)) addrin addrin)))))))))))))))
assign n0001 = sha_state[1:0];
assign n0002 = aes_state[1:0];
assign n0003 = { ( n0001 ), ( n0002 ) };
assign n0004 = 16'h0;
assign n0005 = ( n0003 == n0004 );
assign n0006 = 16'h1;
assign n0007 = ( n0003 == n0006 );
assign n0008 = 16'h2;
assign n0009 = ( n0003 == n0008 );
assign n0010 = 16'h3;
assign n0011 = ( n0003 == n0010 );
assign n0012 = 16'h4;
assign n0013 = ( n0003 == n0012 );
assign n0014 = 16'h5;
assign n0015 = ( n0003 == n0014 );
assign n0016 = 16'h6;
assign n0017 = ( n0003 == n0016 );
assign n0018 = 16'h7;
assign n0019 = ( n0003 == n0018 );
assign n0020 = 16'h8;
assign n0021 = ( n0003 == n0020 );
assign n0022 = 16'h9;
assign n0023 = ( n0003 == n0022 );
assign n0024 = 16'ha;
assign n0025 = ( n0003 == n0024 );
assign n0026 = 16'hb;
assign n0027 = ( n0003 == n0026 );
assign n0028 = 16'hc;
assign n0029 = ( n0003 == n0028 );
assign n0030 = 16'hd;
assign n0031 = ( n0003 == n0030 );
assign n0032 = 16'hf;
assign n0033 = ( aes_bytes_processed + n0032 );
assign n0034 = ( aes_addr + n0033 );
assign n0035 = 16'he;
assign n0036 = ( n0003 == n0035 );
assign n0037 = ( n0036 ) ? ( addrin ) : ( addrin );
assign n0038 = ( n0031 ) ? ( n0034 ) : ( n0037 );
assign n0039 = ( n0029 ) ? ( addrin ) : ( n0038 );
assign n0040 = ( n0027 ) ? ( addrin ) : ( n0039 );
assign n0041 = ( n0025 ) ? ( addrin ) : ( n0040 );
assign n0042 = ( n0023 ) ? ( addrin ) : ( n0041 );
assign n0043 = ( n0021 ) ? ( addrin ) : ( n0042 );
assign n0044 = ( n0019 ) ? ( addrin ) : ( n0043 );
assign n0045 = ( n0017 ) ? ( addrin ) : ( n0044 );
assign n0046 = ( n0015 ) ? ( addrin ) : ( n0045 );
assign n0047 = ( n0013 ) ? ( addrin ) : ( n0046 );
assign n0048 = ( n0011 ) ? ( addrin ) : ( n0047 );
assign n0049 = ( n0009 ) ? ( addrin ) : ( n0048 );
assign n0050 = ( n0007 ) ? ( addrin ) : ( n0049 );
assign n0051 = ( n0005 ) ? ( addrin ) : ( n0050 );
assign RD_xram_0_ADDR = n0051;
// RD_xram_1_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 15 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 63 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 15 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 63 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 63 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 15 16))) (add aes_addr (add aes_bytes_processed (bv 14 16)))))))))
assign n0052 = 16'h3f;
assign n0053 = ( sha_bytes_processed + n0052 );
assign n0054 = ( sha_rdaddr + n0053 );
assign n0055 = ( aes_bytes_processed + n0035 );
assign n0056 = ( aes_addr + n0055 );
assign n0057 = ( n0023 ) ? ( n0034 ) : ( n0056 );
assign n0058 = ( n0019 ) ? ( n0054 ) : ( n0057 );
assign n0059 = ( n0017 ) ? ( n0054 ) : ( n0058 );
assign n0060 = ( n0015 ) ? ( n0034 ) : ( n0059 );
assign n0061 = ( n0013 ) ? ( n0054 ) : ( n0060 );
assign n0062 = ( n0007 ) ? ( n0034 ) : ( n0061 );
assign RD_xram_1_ADDR = n0062;
// RD_xram_2_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 14 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 62 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 14 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 62 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 62 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 14 16))) (add aes_addr (add aes_bytes_processed (bv 13 16)))))))))
assign n0063 = 16'h3e;
assign n0064 = ( sha_bytes_processed + n0063 );
assign n0065 = ( sha_rdaddr + n0064 );
assign n0066 = ( aes_bytes_processed + n0030 );
assign n0067 = ( aes_addr + n0066 );
assign n0068 = ( n0023 ) ? ( n0056 ) : ( n0067 );
assign n0069 = ( n0019 ) ? ( n0065 ) : ( n0068 );
assign n0070 = ( n0017 ) ? ( n0065 ) : ( n0069 );
assign n0071 = ( n0015 ) ? ( n0056 ) : ( n0070 );
assign n0072 = ( n0013 ) ? ( n0065 ) : ( n0071 );
assign n0073 = ( n0007 ) ? ( n0056 ) : ( n0072 );
assign RD_xram_2_ADDR = n0073;
// RD_xram_3_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 13 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 61 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 13 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 61 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 61 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 13 16))) (add aes_addr (add aes_bytes_processed (bv 12 16)))))))))
assign n0074 = 16'h3d;
assign n0075 = ( sha_bytes_processed + n0074 );
assign n0076 = ( sha_rdaddr + n0075 );
assign n0077 = ( aes_bytes_processed + n0028 );
assign n0078 = ( aes_addr + n0077 );
assign n0079 = ( n0023 ) ? ( n0067 ) : ( n0078 );
assign n0080 = ( n0019 ) ? ( n0076 ) : ( n0079 );
assign n0081 = ( n0017 ) ? ( n0076 ) : ( n0080 );
assign n0082 = ( n0015 ) ? ( n0067 ) : ( n0081 );
assign n0083 = ( n0013 ) ? ( n0076 ) : ( n0082 );
assign n0084 = ( n0007 ) ? ( n0067 ) : ( n0083 );
assign RD_xram_3_ADDR = n0084;
// RD_xram_4_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 12 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 60 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 12 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 60 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 60 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 12 16))) (add aes_addr (add aes_bytes_processed (bv 11 16)))))))))
assign n0085 = 16'h3c;
assign n0086 = ( sha_bytes_processed + n0085 );
assign n0087 = ( sha_rdaddr + n0086 );
assign n0088 = ( aes_bytes_processed + n0026 );
assign n0089 = ( aes_addr + n0088 );
assign n0090 = ( n0023 ) ? ( n0078 ) : ( n0089 );
assign n0091 = ( n0019 ) ? ( n0087 ) : ( n0090 );
assign n0092 = ( n0017 ) ? ( n0087 ) : ( n0091 );
assign n0093 = ( n0015 ) ? ( n0078 ) : ( n0092 );
assign n0094 = ( n0013 ) ? ( n0087 ) : ( n0093 );
assign n0095 = ( n0007 ) ? ( n0078 ) : ( n0094 );
assign RD_xram_4_ADDR = n0095;
// RD_xram_5_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 11 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 59 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 11 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 59 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 59 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 11 16))) (add aes_addr (add aes_bytes_processed (bv 10 16)))))))))
assign n0096 = 16'h3b;
assign n0097 = ( sha_bytes_processed + n0096 );
assign n0098 = ( sha_rdaddr + n0097 );
assign n0099 = ( aes_bytes_processed + n0024 );
assign n0100 = ( aes_addr + n0099 );
assign n0101 = ( n0023 ) ? ( n0089 ) : ( n0100 );
assign n0102 = ( n0019 ) ? ( n0098 ) : ( n0101 );
assign n0103 = ( n0017 ) ? ( n0098 ) : ( n0102 );
assign n0104 = ( n0015 ) ? ( n0089 ) : ( n0103 );
assign n0105 = ( n0013 ) ? ( n0098 ) : ( n0104 );
assign n0106 = ( n0007 ) ? ( n0089 ) : ( n0105 );
assign RD_xram_5_ADDR = n0106;
// RD_xram_6_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 10 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 58 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 10 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 58 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 58 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 10 16))) (add aes_addr (add aes_bytes_processed (bv 9 16)))))))))
assign n0107 = 16'h3a;
assign n0108 = ( sha_bytes_processed + n0107 );
assign n0109 = ( sha_rdaddr + n0108 );
assign n0110 = ( aes_bytes_processed + n0022 );
assign n0111 = ( aes_addr + n0110 );
assign n0112 = ( n0023 ) ? ( n0100 ) : ( n0111 );
assign n0113 = ( n0019 ) ? ( n0109 ) : ( n0112 );
assign n0114 = ( n0017 ) ? ( n0109 ) : ( n0113 );
assign n0115 = ( n0015 ) ? ( n0100 ) : ( n0114 );
assign n0116 = ( n0013 ) ? ( n0109 ) : ( n0115 );
assign n0117 = ( n0007 ) ? ( n0100 ) : ( n0116 );
assign RD_xram_6_ADDR = n0117;
// RD_xram_7_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 9 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 57 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 9 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 57 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 57 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 9 16))) (add aes_addr (add aes_bytes_processed (bv 8 16)))))))))
assign n0118 = 16'h39;
assign n0119 = ( sha_bytes_processed + n0118 );
assign n0120 = ( sha_rdaddr + n0119 );
assign n0121 = ( aes_bytes_processed + n0020 );
assign n0122 = ( aes_addr + n0121 );
assign n0123 = ( n0023 ) ? ( n0111 ) : ( n0122 );
assign n0124 = ( n0019 ) ? ( n0120 ) : ( n0123 );
assign n0125 = ( n0017 ) ? ( n0120 ) : ( n0124 );
assign n0126 = ( n0015 ) ? ( n0111 ) : ( n0125 );
assign n0127 = ( n0013 ) ? ( n0120 ) : ( n0126 );
assign n0128 = ( n0007 ) ? ( n0111 ) : ( n0127 );
assign RD_xram_7_ADDR = n0128;
// RD_xram_8_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 8 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 56 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 8 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 56 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 56 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 8 16))) (add aes_addr (add aes_bytes_processed (bv 7 16)))))))))
assign n0129 = 16'h38;
assign n0130 = ( sha_bytes_processed + n0129 );
assign n0131 = ( sha_rdaddr + n0130 );
assign n0132 = ( aes_bytes_processed + n0018 );
assign n0133 = ( aes_addr + n0132 );
assign n0134 = ( n0023 ) ? ( n0122 ) : ( n0133 );
assign n0135 = ( n0019 ) ? ( n0131 ) : ( n0134 );
assign n0136 = ( n0017 ) ? ( n0131 ) : ( n0135 );
assign n0137 = ( n0015 ) ? ( n0122 ) : ( n0136 );
assign n0138 = ( n0013 ) ? ( n0131 ) : ( n0137 );
assign n0139 = ( n0007 ) ? ( n0122 ) : ( n0138 );
assign RD_xram_8_ADDR = n0139;
// RD_xram_9_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 7 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 55 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 7 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 55 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 55 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 7 16))) (add aes_addr (add aes_bytes_processed (bv 6 16)))))))))
assign n0140 = 16'h37;
assign n0141 = ( sha_bytes_processed + n0140 );
assign n0142 = ( sha_rdaddr + n0141 );
assign n0143 = ( aes_bytes_processed + n0016 );
assign n0144 = ( aes_addr + n0143 );
assign n0145 = ( n0023 ) ? ( n0133 ) : ( n0144 );
assign n0146 = ( n0019 ) ? ( n0142 ) : ( n0145 );
assign n0147 = ( n0017 ) ? ( n0142 ) : ( n0146 );
assign n0148 = ( n0015 ) ? ( n0133 ) : ( n0147 );
assign n0149 = ( n0013 ) ? ( n0142 ) : ( n0148 );
assign n0150 = ( n0007 ) ? ( n0133 ) : ( n0149 );
assign RD_xram_9_ADDR = n0150;
// RD_xram_10_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 6 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 54 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 6 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 54 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 54 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 6 16))) (add aes_addr (add aes_bytes_processed (bv 5 16)))))))))
assign n0151 = 16'h36;
assign n0152 = ( sha_bytes_processed + n0151 );
assign n0153 = ( sha_rdaddr + n0152 );
assign n0154 = ( aes_bytes_processed + n0014 );
assign n0155 = ( aes_addr + n0154 );
assign n0156 = ( n0023 ) ? ( n0144 ) : ( n0155 );
assign n0157 = ( n0019 ) ? ( n0153 ) : ( n0156 );
assign n0158 = ( n0017 ) ? ( n0153 ) : ( n0157 );
assign n0159 = ( n0015 ) ? ( n0144 ) : ( n0158 );
assign n0160 = ( n0013 ) ? ( n0153 ) : ( n0159 );
assign n0161 = ( n0007 ) ? ( n0144 ) : ( n0160 );
assign RD_xram_10_ADDR = n0161;
// RD_xram_11_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 5 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 53 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 5 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 53 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 53 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 5 16))) (add aes_addr (add aes_bytes_processed (bv 4 16)))))))))
assign n0162 = 16'h35;
assign n0163 = ( sha_bytes_processed + n0162 );
assign n0164 = ( sha_rdaddr + n0163 );
assign n0165 = ( aes_bytes_processed + n0012 );
assign n0166 = ( aes_addr + n0165 );
assign n0167 = ( n0023 ) ? ( n0155 ) : ( n0166 );
assign n0168 = ( n0019 ) ? ( n0164 ) : ( n0167 );
assign n0169 = ( n0017 ) ? ( n0164 ) : ( n0168 );
assign n0170 = ( n0015 ) ? ( n0155 ) : ( n0169 );
assign n0171 = ( n0013 ) ? ( n0164 ) : ( n0170 );
assign n0172 = ( n0007 ) ? ( n0155 ) : ( n0171 );
assign RD_xram_11_ADDR = n0172;
// RD_xram_12_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 4 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 52 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 4 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 52 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 52 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 4 16))) (add aes_addr (add aes_bytes_processed (bv 3 16)))))))))
assign n0173 = 16'h34;
assign n0174 = ( sha_bytes_processed + n0173 );
assign n0175 = ( sha_rdaddr + n0174 );
assign n0176 = ( aes_bytes_processed + n0010 );
assign n0177 = ( aes_addr + n0176 );
assign n0178 = ( n0023 ) ? ( n0166 ) : ( n0177 );
assign n0179 = ( n0019 ) ? ( n0175 ) : ( n0178 );
assign n0180 = ( n0017 ) ? ( n0175 ) : ( n0179 );
assign n0181 = ( n0015 ) ? ( n0166 ) : ( n0180 );
assign n0182 = ( n0013 ) ? ( n0175 ) : ( n0181 );
assign n0183 = ( n0007 ) ? ( n0166 ) : ( n0182 );
assign RD_xram_12_ADDR = n0183;
// RD_xram_13_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 3 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 51 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 3 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 51 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 51 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 3 16))) (add aes_addr (add aes_bytes_processed (bv 2 16)))))))))
assign n0184 = 16'h33;
assign n0185 = ( sha_bytes_processed + n0184 );
assign n0186 = ( sha_rdaddr + n0185 );
assign n0187 = ( aes_bytes_processed + n0008 );
assign n0188 = ( aes_addr + n0187 );
assign n0189 = ( n0023 ) ? ( n0177 ) : ( n0188 );
assign n0190 = ( n0019 ) ? ( n0186 ) : ( n0189 );
assign n0191 = ( n0017 ) ? ( n0186 ) : ( n0190 );
assign n0192 = ( n0015 ) ? ( n0177 ) : ( n0191 );
assign n0193 = ( n0013 ) ? ( n0186 ) : ( n0192 );
assign n0194 = ( n0007 ) ? ( n0177 ) : ( n0193 );
assign RD_xram_13_ADDR = n0194;
// RD_xram_14_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 2 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 50 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 2 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 50 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 50 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 2 16))) (add aes_addr (add aes_bytes_processed (bv 1 16)))))))))
assign n0195 = 16'h32;
assign n0196 = ( sha_bytes_processed + n0195 );
assign n0197 = ( sha_rdaddr + n0196 );
assign n0198 = ( aes_bytes_processed + n0006 );
assign n0199 = ( aes_addr + n0198 );
assign n0200 = ( n0023 ) ? ( n0188 ) : ( n0199 );
assign n0201 = ( n0019 ) ? ( n0197 ) : ( n0200 );
assign n0202 = ( n0017 ) ? ( n0197 ) : ( n0201 );
assign n0203 = ( n0015 ) ? ( n0188 ) : ( n0202 );
assign n0204 = ( n0013 ) ? ( n0197 ) : ( n0203 );
assign n0205 = ( n0007 ) ? ( n0188 ) : ( n0204 );
assign RD_xram_14_ADDR = n0205;
// RD_xram_15_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 1 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 49 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 1 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 49 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 49 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 1 16))) (add aes_addr (add aes_bytes_processed (bv 0 16)))))))))
assign n0206 = 16'h31;
assign n0207 = ( sha_bytes_processed + n0206 );
assign n0208 = ( sha_rdaddr + n0207 );
assign n0209 = ( aes_bytes_processed + n0004 );
assign n0210 = ( aes_addr + n0209 );
assign n0211 = ( n0023 ) ? ( n0199 ) : ( n0210 );
assign n0212 = ( n0019 ) ? ( n0208 ) : ( n0211 );
assign n0213 = ( n0017 ) ? ( n0208 ) : ( n0212 );
assign n0214 = ( n0015 ) ? ( n0199 ) : ( n0213 );
assign n0215 = ( n0013 ) ? ( n0208 ) : ( n0214 );
assign n0216 = ( n0007 ) ? ( n0199 ) : ( n0215 );
assign RD_xram_15_ADDR = n0216;
// RD_xram_16_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 1 16)) (add aes_addr (add aes_bytes_processed (bv 0 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 48 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add aes_addr (add aes_bytes_processed (bv 0 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 48 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 7 16)) (add sha_rdaddr (add sha_bytes_processed (bv 48 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 9 16)) (add aes_addr (add aes_bytes_processed (bv 0 16))) addrin))))))
assign n0217 = 16'h30;
assign n0218 = ( sha_bytes_processed + n0217 );
assign n0219 = ( sha_rdaddr + n0218 );
assign n0220 = ( n0023 ) ? ( n0210 ) : ( addrin );
assign n0221 = ( n0019 ) ? ( n0219 ) : ( n0220 );
assign n0222 = ( n0017 ) ? ( n0219 ) : ( n0221 );
assign n0223 = ( n0015 ) ? ( n0210 ) : ( n0222 );
assign n0224 = ( n0013 ) ? ( n0219 ) : ( n0223 );
assign n0225 = ( n0007 ) ? ( n0210 ) : ( n0224 );
assign RD_xram_16_ADDR = n0225;
// RD_xram_17_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 47 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 63 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 47 16))) (add sha_rdaddr (add sha_bytes_processed (bv 47 16))))))
assign n0226 = 16'h2f;
assign n0227 = ( sha_bytes_processed + n0226 );
assign n0228 = ( sha_rdaddr + n0227 );
assign n0229 = ( n0017 ) ? ( n0228 ) : ( n0228 );
assign n0230 = ( n0015 ) ? ( n0054 ) : ( n0229 );
assign n0231 = ( n0013 ) ? ( n0228 ) : ( n0230 );
assign RD_xram_17_ADDR = n0231;
// RD_xram_18_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 46 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 62 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 46 16))) (add sha_rdaddr (add sha_bytes_processed (bv 46 16))))))
assign n0232 = 16'h2e;
assign n0233 = ( sha_bytes_processed + n0232 );
assign n0234 = ( sha_rdaddr + n0233 );
assign n0235 = ( n0017 ) ? ( n0234 ) : ( n0234 );
assign n0236 = ( n0015 ) ? ( n0065 ) : ( n0235 );
assign n0237 = ( n0013 ) ? ( n0234 ) : ( n0236 );
assign RD_xram_18_ADDR = n0237;
// RD_xram_19_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 45 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 61 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 45 16))) (add sha_rdaddr (add sha_bytes_processed (bv 45 16))))))
assign n0238 = 16'h2d;
assign n0239 = ( sha_bytes_processed + n0238 );
assign n0240 = ( sha_rdaddr + n0239 );
assign n0241 = ( n0017 ) ? ( n0240 ) : ( n0240 );
assign n0242 = ( n0015 ) ? ( n0076 ) : ( n0241 );
assign n0243 = ( n0013 ) ? ( n0240 ) : ( n0242 );
assign RD_xram_19_ADDR = n0243;
// RD_xram_20_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 44 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 60 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 44 16))) (add sha_rdaddr (add sha_bytes_processed (bv 44 16))))))
assign n0244 = 16'h2c;
assign n0245 = ( sha_bytes_processed + n0244 );
assign n0246 = ( sha_rdaddr + n0245 );
assign n0247 = ( n0017 ) ? ( n0246 ) : ( n0246 );
assign n0248 = ( n0015 ) ? ( n0087 ) : ( n0247 );
assign n0249 = ( n0013 ) ? ( n0246 ) : ( n0248 );
assign RD_xram_20_ADDR = n0249;
// RD_xram_21_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 43 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 59 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 43 16))) (add sha_rdaddr (add sha_bytes_processed (bv 43 16))))))
assign n0250 = 16'h2b;
assign n0251 = ( sha_bytes_processed + n0250 );
assign n0252 = ( sha_rdaddr + n0251 );
assign n0253 = ( n0017 ) ? ( n0252 ) : ( n0252 );
assign n0254 = ( n0015 ) ? ( n0098 ) : ( n0253 );
assign n0255 = ( n0013 ) ? ( n0252 ) : ( n0254 );
assign RD_xram_21_ADDR = n0255;
// RD_xram_22_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 42 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 58 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 42 16))) (add sha_rdaddr (add sha_bytes_processed (bv 42 16))))))
assign n0256 = 16'h2a;
assign n0257 = ( sha_bytes_processed + n0256 );
assign n0258 = ( sha_rdaddr + n0257 );
assign n0259 = ( n0017 ) ? ( n0258 ) : ( n0258 );
assign n0260 = ( n0015 ) ? ( n0109 ) : ( n0259 );
assign n0261 = ( n0013 ) ? ( n0258 ) : ( n0260 );
assign RD_xram_22_ADDR = n0261;
// RD_xram_23_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 41 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 57 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 41 16))) (add sha_rdaddr (add sha_bytes_processed (bv 41 16))))))
assign n0262 = 16'h29;
assign n0263 = ( sha_bytes_processed + n0262 );
assign n0264 = ( sha_rdaddr + n0263 );
assign n0265 = ( n0017 ) ? ( n0264 ) : ( n0264 );
assign n0266 = ( n0015 ) ? ( n0120 ) : ( n0265 );
assign n0267 = ( n0013 ) ? ( n0264 ) : ( n0266 );
assign RD_xram_23_ADDR = n0267;
// RD_xram_24_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 40 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 56 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 40 16))) (add sha_rdaddr (add sha_bytes_processed (bv 40 16))))))
assign n0268 = 16'h28;
assign n0269 = ( sha_bytes_processed + n0268 );
assign n0270 = ( sha_rdaddr + n0269 );
assign n0271 = ( n0017 ) ? ( n0270 ) : ( n0270 );
assign n0272 = ( n0015 ) ? ( n0131 ) : ( n0271 );
assign n0273 = ( n0013 ) ? ( n0270 ) : ( n0272 );
assign RD_xram_24_ADDR = n0273;
// RD_xram_25_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 39 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 55 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 39 16))) (add sha_rdaddr (add sha_bytes_processed (bv 39 16))))))
assign n0274 = 16'h27;
assign n0275 = ( sha_bytes_processed + n0274 );
assign n0276 = ( sha_rdaddr + n0275 );
assign n0277 = ( n0017 ) ? ( n0276 ) : ( n0276 );
assign n0278 = ( n0015 ) ? ( n0142 ) : ( n0277 );
assign n0279 = ( n0013 ) ? ( n0276 ) : ( n0278 );
assign RD_xram_25_ADDR = n0279;
// RD_xram_26_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 38 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 54 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 38 16))) (add sha_rdaddr (add sha_bytes_processed (bv 38 16))))))
assign n0280 = 16'h26;
assign n0281 = ( sha_bytes_processed + n0280 );
assign n0282 = ( sha_rdaddr + n0281 );
assign n0283 = ( n0017 ) ? ( n0282 ) : ( n0282 );
assign n0284 = ( n0015 ) ? ( n0153 ) : ( n0283 );
assign n0285 = ( n0013 ) ? ( n0282 ) : ( n0284 );
assign RD_xram_26_ADDR = n0285;
// RD_xram_27_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 37 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 53 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 37 16))) (add sha_rdaddr (add sha_bytes_processed (bv 37 16))))))
assign n0286 = 16'h25;
assign n0287 = ( sha_bytes_processed + n0286 );
assign n0288 = ( sha_rdaddr + n0287 );
assign n0289 = ( n0017 ) ? ( n0288 ) : ( n0288 );
assign n0290 = ( n0015 ) ? ( n0164 ) : ( n0289 );
assign n0291 = ( n0013 ) ? ( n0288 ) : ( n0290 );
assign RD_xram_27_ADDR = n0291;
// RD_xram_28_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 36 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 52 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 36 16))) (add sha_rdaddr (add sha_bytes_processed (bv 36 16))))))
assign n0292 = 16'h24;
assign n0293 = ( sha_bytes_processed + n0292 );
assign n0294 = ( sha_rdaddr + n0293 );
assign n0295 = ( n0017 ) ? ( n0294 ) : ( n0294 );
assign n0296 = ( n0015 ) ? ( n0175 ) : ( n0295 );
assign n0297 = ( n0013 ) ? ( n0294 ) : ( n0296 );
assign RD_xram_28_ADDR = n0297;
// RD_xram_29_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 35 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 51 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 35 16))) (add sha_rdaddr (add sha_bytes_processed (bv 35 16))))))
assign n0298 = 16'h23;
assign n0299 = ( sha_bytes_processed + n0298 );
assign n0300 = ( sha_rdaddr + n0299 );
assign n0301 = ( n0017 ) ? ( n0300 ) : ( n0300 );
assign n0302 = ( n0015 ) ? ( n0186 ) : ( n0301 );
assign n0303 = ( n0013 ) ? ( n0300 ) : ( n0302 );
assign RD_xram_29_ADDR = n0303;
// RD_xram_30_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 34 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 50 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 34 16))) (add sha_rdaddr (add sha_bytes_processed (bv 34 16))))))
assign n0304 = 16'h22;
assign n0305 = ( sha_bytes_processed + n0304 );
assign n0306 = ( sha_rdaddr + n0305 );
assign n0307 = ( n0017 ) ? ( n0306 ) : ( n0306 );
assign n0308 = ( n0015 ) ? ( n0197 ) : ( n0307 );
assign n0309 = ( n0013 ) ? ( n0306 ) : ( n0308 );
assign RD_xram_30_ADDR = n0309;
// RD_xram_31_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 33 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 49 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 33 16))) (add sha_rdaddr (add sha_bytes_processed (bv 33 16))))))
assign n0310 = 16'h21;
assign n0311 = ( sha_bytes_processed + n0310 );
assign n0312 = ( sha_rdaddr + n0311 );
assign n0313 = ( n0017 ) ? ( n0312 ) : ( n0312 );
assign n0314 = ( n0015 ) ? ( n0208 ) : ( n0313 );
assign n0315 = ( n0013 ) ? ( n0312 ) : ( n0314 );
assign RD_xram_31_ADDR = n0315;
// RD_xram_32_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 32 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 48 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 32 16))) (add sha_rdaddr (add sha_bytes_processed (bv 32 16))))))
assign n0316 = 16'h20;
assign n0317 = ( sha_bytes_processed + n0316 );
assign n0318 = ( sha_rdaddr + n0317 );
assign n0319 = ( n0017 ) ? ( n0318 ) : ( n0318 );
assign n0320 = ( n0015 ) ? ( n0219 ) : ( n0319 );
assign n0321 = ( n0013 ) ? ( n0318 ) : ( n0320 );
assign RD_xram_32_ADDR = n0321;
// RD_xram_33_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 31 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 47 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 31 16))) (add sha_rdaddr (add sha_bytes_processed (bv 31 16))))))
assign n0322 = 16'h1f;
assign n0323 = ( sha_bytes_processed + n0322 );
assign n0324 = ( sha_rdaddr + n0323 );
assign n0325 = ( n0017 ) ? ( n0324 ) : ( n0324 );
assign n0326 = ( n0015 ) ? ( n0228 ) : ( n0325 );
assign n0327 = ( n0013 ) ? ( n0324 ) : ( n0326 );
assign RD_xram_33_ADDR = n0327;
// RD_xram_34_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 30 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 46 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 30 16))) (add sha_rdaddr (add sha_bytes_processed (bv 30 16))))))
assign n0328 = 16'h1e;
assign n0329 = ( sha_bytes_processed + n0328 );
assign n0330 = ( sha_rdaddr + n0329 );
assign n0331 = ( n0017 ) ? ( n0330 ) : ( n0330 );
assign n0332 = ( n0015 ) ? ( n0234 ) : ( n0331 );
assign n0333 = ( n0013 ) ? ( n0330 ) : ( n0332 );
assign RD_xram_34_ADDR = n0333;
// RD_xram_35_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 29 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 45 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 29 16))) (add sha_rdaddr (add sha_bytes_processed (bv 29 16))))))
assign n0334 = 16'h1d;
assign n0335 = ( sha_bytes_processed + n0334 );
assign n0336 = ( sha_rdaddr + n0335 );
assign n0337 = ( n0017 ) ? ( n0336 ) : ( n0336 );
assign n0338 = ( n0015 ) ? ( n0240 ) : ( n0337 );
assign n0339 = ( n0013 ) ? ( n0336 ) : ( n0338 );
assign RD_xram_35_ADDR = n0339;
// RD_xram_36_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 28 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 44 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 28 16))) (add sha_rdaddr (add sha_bytes_processed (bv 28 16))))))
assign n0340 = 16'h1c;
assign n0341 = ( sha_bytes_processed + n0340 );
assign n0342 = ( sha_rdaddr + n0341 );
assign n0343 = ( n0017 ) ? ( n0342 ) : ( n0342 );
assign n0344 = ( n0015 ) ? ( n0246 ) : ( n0343 );
assign n0345 = ( n0013 ) ? ( n0342 ) : ( n0344 );
assign RD_xram_36_ADDR = n0345;
// RD_xram_37_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 27 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 43 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 27 16))) (add sha_rdaddr (add sha_bytes_processed (bv 27 16))))))
assign n0346 = 16'h1b;
assign n0347 = ( sha_bytes_processed + n0346 );
assign n0348 = ( sha_rdaddr + n0347 );
assign n0349 = ( n0017 ) ? ( n0348 ) : ( n0348 );
assign n0350 = ( n0015 ) ? ( n0252 ) : ( n0349 );
assign n0351 = ( n0013 ) ? ( n0348 ) : ( n0350 );
assign RD_xram_37_ADDR = n0351;
// RD_xram_38_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 26 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 42 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 26 16))) (add sha_rdaddr (add sha_bytes_processed (bv 26 16))))))
assign n0352 = 16'h1a;
assign n0353 = ( sha_bytes_processed + n0352 );
assign n0354 = ( sha_rdaddr + n0353 );
assign n0355 = ( n0017 ) ? ( n0354 ) : ( n0354 );
assign n0356 = ( n0015 ) ? ( n0258 ) : ( n0355 );
assign n0357 = ( n0013 ) ? ( n0354 ) : ( n0356 );
assign RD_xram_38_ADDR = n0357;
// RD_xram_39_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 25 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 41 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 25 16))) (add sha_rdaddr (add sha_bytes_processed (bv 25 16))))))
assign n0358 = 16'h19;
assign n0359 = ( sha_bytes_processed + n0358 );
assign n0360 = ( sha_rdaddr + n0359 );
assign n0361 = ( n0017 ) ? ( n0360 ) : ( n0360 );
assign n0362 = ( n0015 ) ? ( n0264 ) : ( n0361 );
assign n0363 = ( n0013 ) ? ( n0360 ) : ( n0362 );
assign RD_xram_39_ADDR = n0363;
// RD_xram_40_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 24 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 40 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 24 16))) (add sha_rdaddr (add sha_bytes_processed (bv 24 16))))))
assign n0364 = 16'h18;
assign n0365 = ( sha_bytes_processed + n0364 );
assign n0366 = ( sha_rdaddr + n0365 );
assign n0367 = ( n0017 ) ? ( n0366 ) : ( n0366 );
assign n0368 = ( n0015 ) ? ( n0270 ) : ( n0367 );
assign n0369 = ( n0013 ) ? ( n0366 ) : ( n0368 );
assign RD_xram_40_ADDR = n0369;
// RD_xram_41_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 23 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 39 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 23 16))) (add sha_rdaddr (add sha_bytes_processed (bv 23 16))))))
assign n0370 = 16'h17;
assign n0371 = ( sha_bytes_processed + n0370 );
assign n0372 = ( sha_rdaddr + n0371 );
assign n0373 = ( n0017 ) ? ( n0372 ) : ( n0372 );
assign n0374 = ( n0015 ) ? ( n0276 ) : ( n0373 );
assign n0375 = ( n0013 ) ? ( n0372 ) : ( n0374 );
assign RD_xram_41_ADDR = n0375;
// RD_xram_42_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 22 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 38 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 22 16))) (add sha_rdaddr (add sha_bytes_processed (bv 22 16))))))
assign n0376 = 16'h16;
assign n0377 = ( sha_bytes_processed + n0376 );
assign n0378 = ( sha_rdaddr + n0377 );
assign n0379 = ( n0017 ) ? ( n0378 ) : ( n0378 );
assign n0380 = ( n0015 ) ? ( n0282 ) : ( n0379 );
assign n0381 = ( n0013 ) ? ( n0378 ) : ( n0380 );
assign RD_xram_42_ADDR = n0381;
// RD_xram_43_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 21 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 37 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 21 16))) (add sha_rdaddr (add sha_bytes_processed (bv 21 16))))))
assign n0382 = 16'h15;
assign n0383 = ( sha_bytes_processed + n0382 );
assign n0384 = ( sha_rdaddr + n0383 );
assign n0385 = ( n0017 ) ? ( n0384 ) : ( n0384 );
assign n0386 = ( n0015 ) ? ( n0288 ) : ( n0385 );
assign n0387 = ( n0013 ) ? ( n0384 ) : ( n0386 );
assign RD_xram_43_ADDR = n0387;
// RD_xram_44_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 20 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 36 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 20 16))) (add sha_rdaddr (add sha_bytes_processed (bv 20 16))))))
assign n0388 = 16'h14;
assign n0389 = ( sha_bytes_processed + n0388 );
assign n0390 = ( sha_rdaddr + n0389 );
assign n0391 = ( n0017 ) ? ( n0390 ) : ( n0390 );
assign n0392 = ( n0015 ) ? ( n0294 ) : ( n0391 );
assign n0393 = ( n0013 ) ? ( n0390 ) : ( n0392 );
assign RD_xram_44_ADDR = n0393;
// RD_xram_45_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 19 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 35 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 19 16))) (add sha_rdaddr (add sha_bytes_processed (bv 19 16))))))
assign n0394 = 16'h13;
assign n0395 = ( sha_bytes_processed + n0394 );
assign n0396 = ( sha_rdaddr + n0395 );
assign n0397 = ( n0017 ) ? ( n0396 ) : ( n0396 );
assign n0398 = ( n0015 ) ? ( n0300 ) : ( n0397 );
assign n0399 = ( n0013 ) ? ( n0396 ) : ( n0398 );
assign RD_xram_45_ADDR = n0399;
// RD_xram_46_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 18 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 34 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 18 16))) (add sha_rdaddr (add sha_bytes_processed (bv 18 16))))))
assign n0400 = 16'h12;
assign n0401 = ( sha_bytes_processed + n0400 );
assign n0402 = ( sha_rdaddr + n0401 );
assign n0403 = ( n0017 ) ? ( n0402 ) : ( n0402 );
assign n0404 = ( n0015 ) ? ( n0306 ) : ( n0403 );
assign n0405 = ( n0013 ) ? ( n0402 ) : ( n0404 );
assign RD_xram_46_ADDR = n0405;
// RD_xram_47_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 17 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 33 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 17 16))) (add sha_rdaddr (add sha_bytes_processed (bv 17 16))))))
assign n0406 = 16'h11;
assign n0407 = ( sha_bytes_processed + n0406 );
assign n0408 = ( sha_rdaddr + n0407 );
assign n0409 = ( n0017 ) ? ( n0408 ) : ( n0408 );
assign n0410 = ( n0015 ) ? ( n0312 ) : ( n0409 );
assign n0411 = ( n0013 ) ? ( n0408 ) : ( n0410 );
assign RD_xram_47_ADDR = n0411;
// RD_xram_48_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 16 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 32 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 16 16))) (add sha_rdaddr (add sha_bytes_processed (bv 16 16))))))
assign n0412 = 16'h10;
assign n0413 = ( sha_bytes_processed + n0412 );
assign n0414 = ( sha_rdaddr + n0413 );
assign n0415 = ( n0017 ) ? ( n0414 ) : ( n0414 );
assign n0416 = ( n0015 ) ? ( n0318 ) : ( n0415 );
assign n0417 = ( n0013 ) ? ( n0414 ) : ( n0416 );
assign RD_xram_48_ADDR = n0417;
// RD_xram_49_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 15 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 31 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 15 16))) (add sha_rdaddr (add sha_bytes_processed (bv 15 16))))))
assign n0418 = ( sha_bytes_processed + n0032 );
assign n0419 = ( sha_rdaddr + n0418 );
assign n0420 = ( n0017 ) ? ( n0419 ) : ( n0419 );
assign n0421 = ( n0015 ) ? ( n0324 ) : ( n0420 );
assign n0422 = ( n0013 ) ? ( n0419 ) : ( n0421 );
assign RD_xram_49_ADDR = n0422;
// RD_xram_50_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 14 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 30 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 14 16))) (add sha_rdaddr (add sha_bytes_processed (bv 14 16))))))
assign n0423 = ( sha_bytes_processed + n0035 );
assign n0424 = ( sha_rdaddr + n0423 );
assign n0425 = ( n0017 ) ? ( n0424 ) : ( n0424 );
assign n0426 = ( n0015 ) ? ( n0330 ) : ( n0425 );
assign n0427 = ( n0013 ) ? ( n0424 ) : ( n0426 );
assign RD_xram_50_ADDR = n0427;
// RD_xram_51_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 13 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 29 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 13 16))) (add sha_rdaddr (add sha_bytes_processed (bv 13 16))))))
assign n0428 = ( sha_bytes_processed + n0030 );
assign n0429 = ( sha_rdaddr + n0428 );
assign n0430 = ( n0017 ) ? ( n0429 ) : ( n0429 );
assign n0431 = ( n0015 ) ? ( n0336 ) : ( n0430 );
assign n0432 = ( n0013 ) ? ( n0429 ) : ( n0431 );
assign RD_xram_51_ADDR = n0432;
// RD_xram_52_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 12 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 28 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 12 16))) (add sha_rdaddr (add sha_bytes_processed (bv 12 16))))))
assign n0433 = ( sha_bytes_processed + n0028 );
assign n0434 = ( sha_rdaddr + n0433 );
assign n0435 = ( n0017 ) ? ( n0434 ) : ( n0434 );
assign n0436 = ( n0015 ) ? ( n0342 ) : ( n0435 );
assign n0437 = ( n0013 ) ? ( n0434 ) : ( n0436 );
assign RD_xram_52_ADDR = n0437;
// RD_xram_53_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 11 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 27 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 11 16))) (add sha_rdaddr (add sha_bytes_processed (bv 11 16))))))
assign n0438 = ( sha_bytes_processed + n0026 );
assign n0439 = ( sha_rdaddr + n0438 );
assign n0440 = ( n0017 ) ? ( n0439 ) : ( n0439 );
assign n0441 = ( n0015 ) ? ( n0348 ) : ( n0440 );
assign n0442 = ( n0013 ) ? ( n0439 ) : ( n0441 );
assign RD_xram_53_ADDR = n0442;
// RD_xram_54_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 10 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 26 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 10 16))) (add sha_rdaddr (add sha_bytes_processed (bv 10 16))))))
assign n0443 = ( sha_bytes_processed + n0024 );
assign n0444 = ( sha_rdaddr + n0443 );
assign n0445 = ( n0017 ) ? ( n0444 ) : ( n0444 );
assign n0446 = ( n0015 ) ? ( n0354 ) : ( n0445 );
assign n0447 = ( n0013 ) ? ( n0444 ) : ( n0446 );
assign RD_xram_54_ADDR = n0447;
// RD_xram_55_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 9 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 25 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 9 16))) (add sha_rdaddr (add sha_bytes_processed (bv 9 16))))))
assign n0448 = ( sha_bytes_processed + n0022 );
assign n0449 = ( sha_rdaddr + n0448 );
assign n0450 = ( n0017 ) ? ( n0449 ) : ( n0449 );
assign n0451 = ( n0015 ) ? ( n0360 ) : ( n0450 );
assign n0452 = ( n0013 ) ? ( n0449 ) : ( n0451 );
assign RD_xram_55_ADDR = n0452;
// RD_xram_56_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 8 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 24 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 8 16))) (add sha_rdaddr (add sha_bytes_processed (bv 8 16))))))
assign n0453 = ( sha_bytes_processed + n0020 );
assign n0454 = ( sha_rdaddr + n0453 );
assign n0455 = ( n0017 ) ? ( n0454 ) : ( n0454 );
assign n0456 = ( n0015 ) ? ( n0366 ) : ( n0455 );
assign n0457 = ( n0013 ) ? ( n0454 ) : ( n0456 );
assign RD_xram_56_ADDR = n0457;
// RD_xram_57_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 7 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 23 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 7 16))) (add sha_rdaddr (add sha_bytes_processed (bv 7 16))))))
assign n0458 = ( sha_bytes_processed + n0018 );
assign n0459 = ( sha_rdaddr + n0458 );
assign n0460 = ( n0017 ) ? ( n0459 ) : ( n0459 );
assign n0461 = ( n0015 ) ? ( n0372 ) : ( n0460 );
assign n0462 = ( n0013 ) ? ( n0459 ) : ( n0461 );
assign RD_xram_57_ADDR = n0462;
// RD_xram_58_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 6 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 22 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 6 16))) (add sha_rdaddr (add sha_bytes_processed (bv 6 16))))))
assign n0463 = ( sha_bytes_processed + n0016 );
assign n0464 = ( sha_rdaddr + n0463 );
assign n0465 = ( n0017 ) ? ( n0464 ) : ( n0464 );
assign n0466 = ( n0015 ) ? ( n0378 ) : ( n0465 );
assign n0467 = ( n0013 ) ? ( n0464 ) : ( n0466 );
assign RD_xram_58_ADDR = n0467;
// RD_xram_59_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 5 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 21 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 5 16))) (add sha_rdaddr (add sha_bytes_processed (bv 5 16))))))
assign n0468 = ( sha_bytes_processed + n0014 );
assign n0469 = ( sha_rdaddr + n0468 );
assign n0470 = ( n0017 ) ? ( n0469 ) : ( n0469 );
assign n0471 = ( n0015 ) ? ( n0384 ) : ( n0470 );
assign n0472 = ( n0013 ) ? ( n0469 ) : ( n0471 );
assign RD_xram_59_ADDR = n0472;
// RD_xram_60_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 4 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 20 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 4 16))) (add sha_rdaddr (add sha_bytes_processed (bv 4 16))))))
assign n0473 = ( sha_bytes_processed + n0012 );
assign n0474 = ( sha_rdaddr + n0473 );
assign n0475 = ( n0017 ) ? ( n0474 ) : ( n0474 );
assign n0476 = ( n0015 ) ? ( n0390 ) : ( n0475 );
assign n0477 = ( n0013 ) ? ( n0474 ) : ( n0476 );
assign RD_xram_60_ADDR = n0477;
// RD_xram_61_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 3 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 19 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 3 16))) (add sha_rdaddr (add sha_bytes_processed (bv 3 16))))))
assign n0478 = ( sha_bytes_processed + n0010 );
assign n0479 = ( sha_rdaddr + n0478 );
assign n0480 = ( n0017 ) ? ( n0479 ) : ( n0479 );
assign n0481 = ( n0015 ) ? ( n0396 ) : ( n0480 );
assign n0482 = ( n0013 ) ? ( n0479 ) : ( n0481 );
assign RD_xram_61_ADDR = n0482;
// RD_xram_62_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 2 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 18 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 2 16))) (add sha_rdaddr (add sha_bytes_processed (bv 2 16))))))
assign n0483 = ( sha_bytes_processed + n0008 );
assign n0484 = ( sha_rdaddr + n0483 );
assign n0485 = ( n0017 ) ? ( n0484 ) : ( n0484 );
assign n0486 = ( n0015 ) ? ( n0402 ) : ( n0485 );
assign n0487 = ( n0013 ) ? ( n0484 ) : ( n0486 );
assign RD_xram_62_ADDR = n0487;
// RD_xram_63_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 1 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 17 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 1 16))) (add sha_rdaddr (add sha_bytes_processed (bv 1 16))))))
assign n0488 = ( sha_bytes_processed + n0006 );
assign n0489 = ( sha_rdaddr + n0488 );
assign n0490 = ( n0017 ) ? ( n0489 ) : ( n0489 );
assign n0491 = ( n0015 ) ? ( n0408 ) : ( n0490 );
assign n0492 = ( n0013 ) ? ( n0489 ) : ( n0491 );
assign RD_xram_63_ADDR = n0492;
// RD_xram_64_ADDR=(if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 4 16)) (add sha_rdaddr (add sha_bytes_processed (bv 0 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 5 16)) (add sha_rdaddr (add sha_bytes_processed (bv 16 16))) (if (eq (concat (extract 1 0 sha_state) (extract 1 0 aes_state)) (bv 6 16)) (add sha_rdaddr (add sha_bytes_processed (bv 0 16))) (add sha_rdaddr (add sha_bytes_processed (bv 0 16))))))
assign n0493 = ( sha_bytes_processed + n0004 );
assign n0494 = ( sha_rdaddr + n0493 );
assign n0495 = ( n0017 ) ? ( n0494 ) : ( n0494 );
assign n0496 = ( n0015 ) ? ( n0414 ) : ( n0495 );
assign n0497 = ( n0013 ) ? ( n0494 ) : ( n0496 );
assign RD_xram_64_ADDR = n0497;
// RD_xram_65_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 15 16)))
assign RD_xram_65_ADDR = n0419;
// RD_xram_66_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 14 16)))
assign RD_xram_66_ADDR = n0424;
// RD_xram_67_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 13 16)))
assign RD_xram_67_ADDR = n0429;
// RD_xram_68_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 12 16)))
assign RD_xram_68_ADDR = n0434;
// RD_xram_69_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 11 16)))
assign RD_xram_69_ADDR = n0439;
// RD_xram_70_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 10 16)))
assign RD_xram_70_ADDR = n0444;
// RD_xram_71_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 9 16)))
assign RD_xram_71_ADDR = n0449;
// RD_xram_72_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 8 16)))
assign RD_xram_72_ADDR = n0454;
// RD_xram_73_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 7 16)))
assign RD_xram_73_ADDR = n0459;
// RD_xram_74_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 6 16)))
assign RD_xram_74_ADDR = n0464;
// RD_xram_75_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 5 16)))
assign RD_xram_75_ADDR = n0469;
// RD_xram_76_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 4 16)))
assign RD_xram_76_ADDR = n0474;
// RD_xram_77_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 3 16)))
assign RD_xram_77_ADDR = n0479;
// RD_xram_78_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 2 16)))
assign RD_xram_78_ADDR = n0484;
// RD_xram_79_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 1 16)))
assign RD_xram_79_ADDR = n0489;
// RD_xram_80_ADDR=(add sha_rdaddr (add sha_bytes_processed (bv 0 16)))
assign RD_xram_80_ADDR = n0494;
// 
// dataout_00
// 
assign n0498 = 16'hff00;
assign n0499 = ( n0498 <= addrin );
assign n0500 = 16'hff40;
assign n0501 = ( addrin < n0500 );
assign n0502 = ( n0499 && n0501 );
assign n0503 = 16'hff06;
assign n0504 = ( n0503 == addrin );
assign n0505 = op[3:2];
assign n0506 = 2'h1;
assign n0507 = ( n0505 == n0506 );
assign n0508 = ( n0504 && n0507 );
assign n0509 = 16'hff02;
assign n0510 = addrin[15:1];
assign n0511 = 1'h0;
assign n0512 = { ( n0510 ), ( n0511 ) };
assign n0513 = ( n0509 == n0512 );
assign n0514 = ( n0513 && n0507 );
assign n0515 = addrin[0:0];
assign n0516 = ( n0515 == n0511 );
assign n0517 = aes_addr[7:0];
assign n0518 = aes_addr[15:8];
assign n0519 = ( n0516 ) ? ( n0517 ) : ( n0518 );
assign n0520 = 16'hff04;
assign n0521 = ( n0520 == n0512 );
assign n0522 = ( n0521 && n0507 );
assign n0523 = aes_len[7:0];
assign n0524 = aes_len[15:8];
assign n0525 = ( n0516 ) ? ( n0523 ) : ( n0524 );
assign n0526 = 16'hff10;
assign n0527 = addrin[15:4];
assign n0528 = 4'h0;
assign n0529 = { ( n0527 ), ( n0528 ) };
assign n0530 = ( n0526 == n0529 );
assign n0531 = ( n0530 && n0507 );
assign n0532 = addrin[3:0];
assign n0533 = ( n0532 == n0528 );
assign n0534 = aes_ctr[7:0];
assign n0535 = 4'h1;
assign n0536 = ( n0532 == n0535 );
assign n0537 = aes_ctr[15:8];
assign n0538 = 4'h2;
assign n0539 = ( n0532 == n0538 );
assign n0540 = aes_ctr[23:16];
assign n0541 = 4'h3;
assign n0542 = ( n0532 == n0541 );
assign n0543 = aes_ctr[31:24];
assign n0544 = 4'h4;
assign n0545 = ( n0532 == n0544 );
assign n0546 = aes_ctr[39:32];
assign n0547 = 4'h5;
assign n0548 = ( n0532 == n0547 );
assign n0549 = aes_ctr[47:40];
assign n0550 = 4'h6;
assign n0551 = ( n0532 == n0550 );
assign n0552 = aes_ctr[55:48];
assign n0553 = 4'h7;
assign n0554 = ( n0532 == n0553 );
assign n0555 = aes_ctr[63:56];
assign n0556 = 4'h8;
assign n0557 = ( n0532 == n0556 );
assign n0558 = aes_ctr[71:64];
assign n0559 = 4'h9;
assign n0560 = ( n0532 == n0559 );
assign n0561 = aes_ctr[79:72];
assign n0562 = 4'ha;
assign n0563 = ( n0532 == n0562 );
assign n0564 = aes_ctr[87:80];
assign n0565 = 4'hb;
assign n0566 = ( n0532 == n0565 );
assign n0567 = aes_ctr[95:88];
assign n0568 = 4'hc;
assign n0569 = ( n0532 == n0568 );
assign n0570 = aes_ctr[103:96];
assign n0571 = 4'hd;
assign n0572 = ( n0532 == n0571 );
assign n0573 = aes_ctr[111:104];
assign n0574 = 4'he;
assign n0575 = ( n0532 == n0574 );
assign n0576 = aes_ctr[119:112];
assign n0577 = aes_ctr[127:120];
assign n0578 = ( n0575 ) ? ( n0576 ) : ( n0577 );
assign n0579 = ( n0572 ) ? ( n0573 ) : ( n0578 );
assign n0580 = ( n0569 ) ? ( n0570 ) : ( n0579 );
assign n0581 = ( n0566 ) ? ( n0567 ) : ( n0580 );
assign n0582 = ( n0563 ) ? ( n0564 ) : ( n0581 );
assign n0583 = ( n0560 ) ? ( n0561 ) : ( n0582 );
assign n0584 = ( n0557 ) ? ( n0558 ) : ( n0583 );
assign n0585 = ( n0554 ) ? ( n0555 ) : ( n0584 );
assign n0586 = ( n0551 ) ? ( n0552 ) : ( n0585 );
assign n0587 = ( n0548 ) ? ( n0549 ) : ( n0586 );
assign n0588 = ( n0545 ) ? ( n0546 ) : ( n0587 );
assign n0589 = ( n0542 ) ? ( n0543 ) : ( n0588 );
assign n0590 = ( n0539 ) ? ( n0540 ) : ( n0589 );
assign n0591 = ( n0536 ) ? ( n0537 ) : ( n0590 );
assign n0592 = ( n0533 ) ? ( n0534 ) : ( n0591 );
assign n0593 = 16'hff20;
assign n0594 = ( n0593 == n0529 );
assign n0595 = ( n0594 && n0507 );
assign n0596 = aes_key0[7:0];
assign n0597 = aes_key0[15:8];
assign n0598 = aes_key0[23:16];
assign n0599 = aes_key0[31:24];
assign n0600 = aes_key0[39:32];
assign n0601 = aes_key0[47:40];
assign n0602 = aes_key0[55:48];
assign n0603 = aes_key0[63:56];
assign n0604 = aes_key0[71:64];
assign n0605 = aes_key0[79:72];
assign n0606 = aes_key0[87:80];
assign n0607 = aes_key0[95:88];
assign n0608 = aes_key0[103:96];
assign n0609 = aes_key0[111:104];
assign n0610 = aes_key0[119:112];
assign n0611 = aes_key0[127:120];
assign n0612 = ( n0575 ) ? ( n0610 ) : ( n0611 );
assign n0613 = ( n0572 ) ? ( n0609 ) : ( n0612 );
assign n0614 = ( n0569 ) ? ( n0608 ) : ( n0613 );
assign n0615 = ( n0566 ) ? ( n0607 ) : ( n0614 );
assign n0616 = ( n0563 ) ? ( n0606 ) : ( n0615 );
assign n0617 = ( n0560 ) ? ( n0605 ) : ( n0616 );
assign n0618 = ( n0557 ) ? ( n0604 ) : ( n0617 );
assign n0619 = ( n0554 ) ? ( n0603 ) : ( n0618 );
assign n0620 = ( n0551 ) ? ( n0602 ) : ( n0619 );
assign n0621 = ( n0548 ) ? ( n0601 ) : ( n0620 );
assign n0622 = ( n0545 ) ? ( n0600 ) : ( n0621 );
assign n0623 = ( n0542 ) ? ( n0599 ) : ( n0622 );
assign n0624 = ( n0539 ) ? ( n0598 ) : ( n0623 );
assign n0625 = ( n0536 ) ? ( n0597 ) : ( n0624 );
assign n0626 = ( n0533 ) ? ( n0596 ) : ( n0625 );
assign n0627 = 16'hff30;
assign n0628 = ( n0627 == n0529 );
assign n0629 = ( n0628 && n0507 );
assign n0630 = aes_key1[7:0];
assign n0631 = aes_key1[15:8];
assign n0632 = aes_key1[23:16];
assign n0633 = aes_key1[31:24];
assign n0634 = aes_key1[39:32];
assign n0635 = aes_key1[47:40];
assign n0636 = aes_key1[55:48];
assign n0637 = aes_key1[63:56];
assign n0638 = aes_key1[71:64];
assign n0639 = aes_key1[79:72];
assign n0640 = aes_key1[87:80];
assign n0641 = aes_key1[95:88];
assign n0642 = aes_key1[103:96];
assign n0643 = aes_key1[111:104];
assign n0644 = aes_key1[119:112];
assign n0645 = aes_key1[127:120];
assign n0646 = ( n0575 ) ? ( n0644 ) : ( n0645 );
assign n0647 = ( n0572 ) ? ( n0643 ) : ( n0646 );
assign n0648 = ( n0569 ) ? ( n0642 ) : ( n0647 );
assign n0649 = ( n0566 ) ? ( n0641 ) : ( n0648 );
assign n0650 = ( n0563 ) ? ( n0640 ) : ( n0649 );
assign n0651 = ( n0560 ) ? ( n0639 ) : ( n0650 );
assign n0652 = ( n0557 ) ? ( n0638 ) : ( n0651 );
assign n0653 = ( n0554 ) ? ( n0637 ) : ( n0652 );
assign n0654 = ( n0551 ) ? ( n0636 ) : ( n0653 );
assign n0655 = ( n0548 ) ? ( n0635 ) : ( n0654 );
assign n0656 = ( n0545 ) ? ( n0634 ) : ( n0655 );
assign n0657 = ( n0542 ) ? ( n0633 ) : ( n0656 );
assign n0658 = ( n0539 ) ? ( n0632 ) : ( n0657 );
assign n0659 = ( n0536 ) ? ( n0631 ) : ( n0658 );
assign n0660 = ( n0533 ) ? ( n0630 ) : ( n0659 );
assign n0661 = 8'h0;
assign n0662 = ( n0629 ) ? ( n0660 ) : ( n0661 );
assign n0663 = ( n0595 ) ? ( n0626 ) : ( n0662 );
assign n0664 = ( n0531 ) ? ( n0592 ) : ( n0663 );
assign n0665 = ( n0522 ) ? ( n0525 ) : ( n0664 );
assign n0666 = ( n0514 ) ? ( n0519 ) : ( n0665 );
assign n0667 = ( n0508 ) ? ( aes_state ) : ( n0666 );
assign n0668 = 16'hfe00;
assign n0669 = ( n0668 <= addrin );
assign n0670 = 16'hfe10;
assign n0671 = ( addrin < n0670 );
assign n0672 = ( n0669 && n0671 );
assign n0673 = ( n0668 == addrin );
assign n0674 = ( n0673 && n0507 );
assign n0675 = 16'hfe02;
assign n0676 = ( n0675 == n0512 );
assign n0677 = ( n0676 && n0507 );
assign n0678 = sha_rdaddr[7:0];
assign n0679 = sha_rdaddr[15:8];
assign n0680 = ( n0516 ) ? ( n0678 ) : ( n0679 );
assign n0681 = 16'hfe04;
assign n0682 = ( n0681 == n0512 );
assign n0683 = ( n0682 && n0507 );
assign n0684 = sha_wraddr[7:0];
assign n0685 = sha_wraddr[15:8];
assign n0686 = ( n0516 ) ? ( n0684 ) : ( n0685 );
assign n0687 = 16'hfe06;
assign n0688 = ( n0687 == n0512 );
assign n0689 = ( n0688 && n0507 );
assign n0690 = sha_len[7:0];
assign n0691 = sha_len[15:8];
assign n0692 = ( n0516 ) ? ( n0690 ) : ( n0691 );
assign n0693 = ( n0689 ) ? ( n0692 ) : ( n0661 );
assign n0694 = ( n0683 ) ? ( n0686 ) : ( n0693 );
assign n0695 = ( n0677 ) ? ( n0680 ) : ( n0694 );
assign n0696 = ( n0674 ) ? ( sha_state ) : ( n0695 );
assign n0697 = ( n0507 ) ? ( RD_xram_0 ) : ( n0661 );
assign n0698 = ( n0672 ) ? ( n0696 ) : ( n0697 );
assign n0699 = ( n0502 ) ? ( n0667 ) : ( n0698 );
assign dataout_00 = n0699;
// 
// sha_rdaddr_00
// 
assign n0700 = 2'h2;
assign n0701 = ( n0505 == n0700 );
assign n0702 = ( n0676 && n0701 );
assign n0703 = { ( n0679 ), ( datain ) };
assign n0704 = { ( datain ), ( n0678 ) };
assign n0705 = ( n0516 ) ? ( n0703 ) : ( n0704 );
assign n0706 = ( n0702 ) ? ( n0705 ) : ( sha_rdaddr );
assign sha_rdaddr_00 = n0706;
// 
// aes_addr_00
// 
assign n0707 = ( aes_state == n0661 );
assign n0708 = ( n0701 && n0707 );
assign n0709 = ( n0513 && n0708 );
assign n0710 = { ( n0518 ), ( datain ) };
assign n0711 = { ( datain ), ( n0517 ) };
assign n0712 = ( n0516 ) ? ( n0710 ) : ( n0711 );
assign n0713 = ( n0709 ) ? ( n0712 ) : ( aes_addr );
assign aes_addr_00 = n0713;
// 
// aes_ctr_00
// 
assign n0714 = ( n0530 && n0708 );
assign n0715 = aes_ctr[127:8];
assign n0716 = { ( n0715 ), ( datain ) };
assign n0717 = aes_ctr[127:16];
assign n0718 = { ( n0717 ), ( datain ), ( n0534 ) };
assign n0719 = aes_ctr[127:24];
assign n0720 = aes_ctr[15:0];
assign n0721 = { ( n0719 ), ( datain ), ( n0720 ) };
assign n0722 = aes_ctr[127:32];
assign n0723 = aes_ctr[23:0];
assign n0724 = { ( n0722 ), ( datain ), ( n0723 ) };
assign n0725 = aes_ctr[127:40];
assign n0726 = aes_ctr[31:0];
assign n0727 = { ( n0725 ), ( datain ), ( n0726 ) };
assign n0728 = aes_ctr[127:48];
assign n0729 = aes_ctr[39:0];
assign n0730 = { ( n0728 ), ( datain ), ( n0729 ) };
assign n0731 = aes_ctr[127:56];
assign n0732 = aes_ctr[47:0];
assign n0733 = { ( n0731 ), ( datain ), ( n0732 ) };
assign n0734 = aes_ctr[127:64];
assign n0735 = aes_ctr[55:0];
assign n0736 = { ( n0734 ), ( datain ), ( n0735 ) };
assign n0737 = aes_ctr[127:72];
assign n0738 = aes_ctr[63:0];
assign n0739 = { ( n0737 ), ( datain ), ( n0738 ) };
assign n0740 = aes_ctr[127:80];
assign n0741 = aes_ctr[71:0];
assign n0742 = { ( n0740 ), ( datain ), ( n0741 ) };
assign n0743 = aes_ctr[127:88];
assign n0744 = aes_ctr[79:0];
assign n0745 = { ( n0743 ), ( datain ), ( n0744 ) };
assign n0746 = aes_ctr[127:96];
assign n0747 = aes_ctr[87:0];
assign n0748 = { ( n0746 ), ( datain ), ( n0747 ) };
assign n0749 = aes_ctr[127:104];
assign n0750 = aes_ctr[95:0];
assign n0751 = { ( n0749 ), ( datain ), ( n0750 ) };
assign n0752 = aes_ctr[127:112];
assign n0753 = aes_ctr[103:0];
assign n0754 = { ( n0752 ), ( datain ), ( n0753 ) };
assign n0755 = aes_ctr[111:0];
assign n0756 = { ( n0577 ), ( datain ), ( n0755 ) };
assign n0757 = aes_ctr[119:0];
assign n0758 = { ( datain ), ( n0757 ) };
assign n0759 = ( n0575 ) ? ( n0756 ) : ( n0758 );
assign n0760 = ( n0572 ) ? ( n0754 ) : ( n0759 );
assign n0761 = ( n0569 ) ? ( n0751 ) : ( n0760 );
assign n0762 = ( n0566 ) ? ( n0748 ) : ( n0761 );
assign n0763 = ( n0563 ) ? ( n0745 ) : ( n0762 );
assign n0764 = ( n0560 ) ? ( n0742 ) : ( n0763 );
assign n0765 = ( n0557 ) ? ( n0739 ) : ( n0764 );
assign n0766 = ( n0554 ) ? ( n0736 ) : ( n0765 );
assign n0767 = ( n0551 ) ? ( n0733 ) : ( n0766 );
assign n0768 = ( n0548 ) ? ( n0730 ) : ( n0767 );
assign n0769 = ( n0545 ) ? ( n0727 ) : ( n0768 );
assign n0770 = ( n0542 ) ? ( n0724 ) : ( n0769 );
assign n0771 = ( n0539 ) ? ( n0721 ) : ( n0770 );
assign n0772 = ( n0536 ) ? ( n0718 ) : ( n0771 );
assign n0773 = ( n0533 ) ? ( n0716 ) : ( n0772 );
assign n0774 = ( n0714 ) ? ( n0773 ) : ( aes_ctr );
assign aes_ctr_00 = n0774;
// 
// aes_bytes_processed_00
// 
assign n0775 = datain[0:0];
assign n0776 = 1'h1;
assign n0777 = ( n0775 == n0776 );
assign n0778 = ( n0498 == addrin );
assign n0779 = ( n0777 && n0708 && n0778 );
assign n0780 = ( n0779 ) ? ( n0004 ) : ( aes_bytes_processed );
assign aes_bytes_processed_00 = n0780;
// 
// sha_len_00
// 
assign n0781 = ( n0688 && n0701 );
assign n0782 = { ( n0691 ), ( datain ) };
assign n0783 = { ( datain ), ( n0690 ) };
assign n0784 = ( n0516 ) ? ( n0782 ) : ( n0783 );
assign n0785 = ( n0781 ) ? ( n0784 ) : ( sha_len );
assign sha_len_00 = n0785;
// 
// aes_key1_00
// 
assign n0786 = ( n0628 && n0708 );
assign n0787 = aes_key1[127:8];
assign n0788 = { ( n0787 ), ( datain ) };
assign n0789 = aes_key1[127:16];
assign n0790 = { ( n0789 ), ( datain ), ( n0630 ) };
assign n0791 = aes_key1[127:24];
assign n0792 = aes_key1[15:0];
assign n0793 = { ( n0791 ), ( datain ), ( n0792 ) };
assign n0794 = aes_key1[127:32];
assign n0795 = aes_key1[23:0];
assign n0796 = { ( n0794 ), ( datain ), ( n0795 ) };
assign n0797 = aes_key1[127:40];
assign n0798 = aes_key1[31:0];
assign n0799 = { ( n0797 ), ( datain ), ( n0798 ) };
assign n0800 = aes_key1[127:48];
assign n0801 = aes_key1[39:0];
assign n0802 = { ( n0800 ), ( datain ), ( n0801 ) };
assign n0803 = aes_key1[127:56];
assign n0804 = aes_key1[47:0];
assign n0805 = { ( n0803 ), ( datain ), ( n0804 ) };
assign n0806 = aes_key1[127:64];
assign n0807 = aes_key1[55:0];
assign n0808 = { ( n0806 ), ( datain ), ( n0807 ) };
assign n0809 = aes_key1[127:72];
assign n0810 = aes_key1[63:0];
assign n0811 = { ( n0809 ), ( datain ), ( n0810 ) };
assign n0812 = aes_key1[127:80];
assign n0813 = aes_key1[71:0];
assign n0814 = { ( n0812 ), ( datain ), ( n0813 ) };
assign n0815 = aes_key1[127:88];
assign n0816 = aes_key1[79:0];
assign n0817 = { ( n0815 ), ( datain ), ( n0816 ) };
assign n0818 = aes_key1[127:96];
assign n0819 = aes_key1[87:0];
assign n0820 = { ( n0818 ), ( datain ), ( n0819 ) };
assign n0821 = aes_key1[127:104];
assign n0822 = aes_key1[95:0];
assign n0823 = { ( n0821 ), ( datain ), ( n0822 ) };
assign n0824 = aes_key1[127:112];
assign n0825 = aes_key1[103:0];
assign n0826 = { ( n0824 ), ( datain ), ( n0825 ) };
assign n0827 = aes_key1[111:0];
assign n0828 = { ( n0645 ), ( datain ), ( n0827 ) };
assign n0829 = aes_key1[119:0];
assign n0830 = { ( datain ), ( n0829 ) };
assign n0831 = ( n0575 ) ? ( n0828 ) : ( n0830 );
assign n0832 = ( n0572 ) ? ( n0826 ) : ( n0831 );
assign n0833 = ( n0569 ) ? ( n0823 ) : ( n0832 );
assign n0834 = ( n0566 ) ? ( n0820 ) : ( n0833 );
assign n0835 = ( n0563 ) ? ( n0817 ) : ( n0834 );
assign n0836 = ( n0560 ) ? ( n0814 ) : ( n0835 );
assign n0837 = ( n0557 ) ? ( n0811 ) : ( n0836 );
assign n0838 = ( n0554 ) ? ( n0808 ) : ( n0837 );
assign n0839 = ( n0551 ) ? ( n0805 ) : ( n0838 );
assign n0840 = ( n0548 ) ? ( n0802 ) : ( n0839 );
assign n0841 = ( n0545 ) ? ( n0799 ) : ( n0840 );
assign n0842 = ( n0542 ) ? ( n0796 ) : ( n0841 );
assign n0843 = ( n0539 ) ? ( n0793 ) : ( n0842 );
assign n0844 = ( n0536 ) ? ( n0790 ) : ( n0843 );
assign n0845 = ( n0533 ) ? ( n0788 ) : ( n0844 );
assign n0846 = ( n0786 ) ? ( n0845 ) : ( aes_key1 );
assign aes_key1_00 = n0846;
// 
// aes_key0_00
// 
assign n0847 = ( n0594 && n0708 );
assign n0848 = aes_key0[127:8];
assign n0849 = { ( n0848 ), ( datain ) };
assign n0850 = aes_key0[127:16];
assign n0851 = { ( n0850 ), ( datain ), ( n0596 ) };
assign n0852 = aes_key0[127:24];
assign n0853 = aes_key0[15:0];
assign n0854 = { ( n0852 ), ( datain ), ( n0853 ) };
assign n0855 = aes_key0[127:32];
assign n0856 = aes_key0[23:0];
assign n0857 = { ( n0855 ), ( datain ), ( n0856 ) };
assign n0858 = aes_key0[127:40];
assign n0859 = aes_key0[31:0];
assign n0860 = { ( n0858 ), ( datain ), ( n0859 ) };
assign n0861 = aes_key0[127:48];
assign n0862 = aes_key0[39:0];
assign n0863 = { ( n0861 ), ( datain ), ( n0862 ) };
assign n0864 = aes_key0[127:56];
assign n0865 = aes_key0[47:0];
assign n0866 = { ( n0864 ), ( datain ), ( n0865 ) };
assign n0867 = aes_key0[127:64];
assign n0868 = aes_key0[55:0];
assign n0869 = { ( n0867 ), ( datain ), ( n0868 ) };
assign n0870 = aes_key0[127:72];
assign n0871 = aes_key0[63:0];
assign n0872 = { ( n0870 ), ( datain ), ( n0871 ) };
assign n0873 = aes_key0[127:80];
assign n0874 = aes_key0[71:0];
assign n0875 = { ( n0873 ), ( datain ), ( n0874 ) };
assign n0876 = aes_key0[127:88];
assign n0877 = aes_key0[79:0];
assign n0878 = { ( n0876 ), ( datain ), ( n0877 ) };
assign n0879 = aes_key0[127:96];
assign n0880 = aes_key0[87:0];
assign n0881 = { ( n0879 ), ( datain ), ( n0880 ) };
assign n0882 = aes_key0[127:104];
assign n0883 = aes_key0[95:0];
assign n0884 = { ( n0882 ), ( datain ), ( n0883 ) };
assign n0885 = aes_key0[127:112];
assign n0886 = aes_key0[103:0];
assign n0887 = { ( n0885 ), ( datain ), ( n0886 ) };
assign n0888 = aes_key0[111:0];
assign n0889 = { ( n0611 ), ( datain ), ( n0888 ) };
assign n0890 = aes_key0[119:0];
assign n0891 = { ( datain ), ( n0890 ) };
assign n0892 = ( n0575 ) ? ( n0889 ) : ( n0891 );
assign n0893 = ( n0572 ) ? ( n0887 ) : ( n0892 );
assign n0894 = ( n0569 ) ? ( n0884 ) : ( n0893 );
assign n0895 = ( n0566 ) ? ( n0881 ) : ( n0894 );
assign n0896 = ( n0563 ) ? ( n0878 ) : ( n0895 );
assign n0897 = ( n0560 ) ? ( n0875 ) : ( n0896 );
assign n0898 = ( n0557 ) ? ( n0872 ) : ( n0897 );
assign n0899 = ( n0554 ) ? ( n0869 ) : ( n0898 );
assign n0900 = ( n0551 ) ? ( n0866 ) : ( n0899 );
assign n0901 = ( n0548 ) ? ( n0863 ) : ( n0900 );
assign n0902 = ( n0545 ) ? ( n0860 ) : ( n0901 );
assign n0903 = ( n0542 ) ? ( n0857 ) : ( n0902 );
assign n0904 = ( n0539 ) ? ( n0854 ) : ( n0903 );
assign n0905 = ( n0536 ) ? ( n0851 ) : ( n0904 );
assign n0906 = ( n0533 ) ? ( n0849 ) : ( n0905 );
assign n0907 = ( n0847 ) ? ( n0906 ) : ( aes_key0 );
assign aes_key0_00 = n0907;
// 
// aes_len_00
// 
assign n0908 = ( n0521 && n0708 );
assign n0909 = { ( n0524 ), ( datain ) };
assign n0910 = { ( datain ), ( n0523 ) };
assign n0911 = ( n0516 ) ? ( n0909 ) : ( n0910 );
assign n0912 = ( n0908 ) ? ( n0911 ) : ( aes_len );
assign aes_len_00 = n0912;
// 
// sha_state_00
// 
assign n0913 = ( sha_state == n0661 );
assign n0914 = ( n0701 && n0913 );
assign n0915 = ( n0777 && n0914 && n0673 );
assign n0916 = 8'h1;
assign n0917 = ( n0915 ) ? ( n0916 ) : ( n0661 );
assign sha_state_00 = n0917;
// 
// sha_bytes_processed_00
// 
assign n0918 = ( n0915 ) ? ( n0004 ) : ( sha_bytes_processed );
assign sha_bytes_processed_00 = n0918;
// 
// sha_wraddr_00
// 
assign n0919 = ( n0682 && n0701 );
assign n0920 = { ( n0685 ), ( datain ) };
assign n0921 = { ( datain ), ( n0684 ) };
assign n0922 = ( n0516 ) ? ( n0920 ) : ( n0921 );
assign n0923 = ( n0919 ) ? ( n0922 ) : ( sha_wraddr );
assign sha_wraddr_00 = n0923;
// 
// sha_digest_00
// 
assign n0924 = ( sha_state == n0916 );
assign n0925 = 160'h0;
assign n0926 = ( n0915 ) ? ( n0925 ) : ( sha_digest );
assign n0927 = 8'h2;
assign n0928 = ( sha_state == n0927 );
assign n0929 = op[1:1];
assign n0930 = ( n0929 == n0776 );
assign n0931 = { ( input_sha_func_0 ), ( input_sha_func_1 ), ( input_sha_func_2 ) };
assign n0932 = ( n0930 ) ? ( n0931 ) : ( sha_digest );
assign n0933 = ( n0928 ) ? ( n0932 ) : ( sha_digest );
assign n0934 = ( n0924 ) ? ( n0926 ) : ( n0933 );
assign sha_digest_00 = n0934;
// 
// xram_00
// 
// 
// aes_state_00
// 
assign n0935 = ( n0779 ) ? ( n0916 ) : ( n0661 );
assign aes_state_00 = n0935;
assign n0936 = !( n0502 );
assign n0937 = !( n0672 );
assign n0938 = ( n0701 && n0936 && n0937 );
assign n0939 = ( 1 && n0938 );
assign WR_XRAM_EN_00 = n0939;
assign WR_XRAM_ADDR_00 = addrin;
// 
// dataout_01
// 
assign n0940 = 16'hff01;
assign n0941 = ( n0940 == addrin );
assign n0942 = ( n0941 && n0507 );
assign n0943 = ( n0942 ) ? ( aes_state ) : ( n0666 );
assign n0944 = 16'hfe0c;
assign n0945 = ( n0944 == addrin );
assign n0946 = ( n0945 && n0507 );
assign n0947 = ( n0946 ) ? ( sha_state ) : ( n0695 );
assign n0948 = ( n0672 ) ? ( n0947 ) : ( n0697 );
assign n0949 = ( n0502 ) ? ( n0943 ) : ( n0948 );
assign dataout_01 = n0949;
// 
// sha_rdaddr_01
// 
assign sha_rdaddr_01 = n0706;
// 
// aes_bytes_processed_01
// 
assign n0950 = 16'hff38;
assign n0951 = ( n0950 == addrin );
assign n0952 = ( n0777 && n0708 && n0951 );
assign n0953 = ( n0952 ) ? ( n0004 ) : ( aes_bytes_processed );
assign aes_bytes_processed_01 = n0953;
// 
// sha_len_01
// 
assign sha_len_01 = n0785;
// 
// aes_read_data_01
// 
assign n0954 = op[0:0];
assign n0955 = ( n0954 == n0776 );
assign n0956 = { ( RD_xram_1 ), ( RD_xram_2 ), ( RD_xram_3 ), ( RD_xram_4 ), ( RD_xram_5 ), ( RD_xram_6 ), ( RD_xram_7 ), ( RD_xram_8 ), ( RD_xram_9 ), ( RD_xram_10 ), ( RD_xram_11 ), ( RD_xram_12 ), ( RD_xram_13 ), ( RD_xram_14 ), ( RD_xram_15 ), ( RD_xram_16 ) };
assign n0957 = ( n0955 ) ? ( n0956 ) : ( aes_read_data );
assign aes_read_data_01 = n0957;
// 
// sha_bytes_processed_01
// 
assign sha_bytes_processed_01 = n0918;
// 
// sha_wraddr_01
// 
assign sha_wraddr_01 = n0923;
// 
// sha_digest_01
// 
assign n0958 = { ( input_sha_func_3 ), ( input_sha_func_4 ), ( input_sha_func_5 ) };
assign n0959 = ( n0930 ) ? ( n0958 ) : ( sha_digest );
assign n0960 = ( n0928 ) ? ( n0959 ) : ( sha_digest );
assign n0961 = ( n0924 ) ? ( n0926 ) : ( n0960 );
assign sha_digest_01 = n0961;
// 
// xram_01
// 
// 
// aes_state_01
// 
assign n0962 = ( n0955 ) ? ( n0927 ) : ( n0916 );
assign aes_state_01 = n0962;
// 
// sha_state_01
// 
assign sha_state_01 = n0917;
assign WR_XRAM_EN_01 = n0939;
assign WR_XRAM_ADDR_01 = addrin;
// 
// sha_rdaddr_02
// 
assign sha_rdaddr_02 = n0706;
// 
// aes_bytes_processed_02
// 
assign aes_bytes_processed_02 = n0953;
// 
// sha_len_02
// 
assign sha_len_02 = n0785;
// 
// sha_state_02
// 
assign sha_state_02 = n0917;
// 
// sha_bytes_processed_02
// 
assign sha_bytes_processed_02 = n0918;
// 
// sha_wraddr_02
// 
assign sha_wraddr_02 = n0923;
// 
// dataout_02
// 
assign n0963 = ( n0502 ) ? ( n0943 ) : ( n0698 );
assign dataout_02 = n0963;
// 
// xram_02
// 
// 
// aes_state_02
// 
assign n0964 = 8'h3;
assign n0965 = ( n0955 ) ? ( n0964 ) : ( n0927 );
assign aes_state_02 = n0965;
// 
// aes_enc_data_02
// 
assign n0966 = { ( input_aes_func_6 ), ( input_aes_func_7 ) };
assign n0967 = ( n0955 ) ? ( n0966 ) : ( aes_enc_data );
assign aes_enc_data_02 = n0967;
// 
// sha_digest_02
// 
assign n0968 = { ( input_sha_func_8 ), ( input_sha_func_9 ), ( input_sha_func_10 ) };
assign n0969 = ( n0930 ) ? ( n0968 ) : ( sha_digest );
assign n0970 = ( n0928 ) ? ( n0969 ) : ( sha_digest );
assign n0971 = ( n0924 ) ? ( n0926 ) : ( n0970 );
assign sha_digest_02 = n0971;
assign WR_XRAM_EN_02 = n0939;
assign WR_XRAM_ADDR_02 = addrin;
// 
// xram_03
// 
// 
// aes_bytes_processed_03
// 
assign n0972 = ( aes_bytes_processed + n0412 );
assign n0973 = ( n0955 ) ? ( n0972 ) : ( aes_bytes_processed );
assign aes_bytes_processed_03 = n0973;
// 
// sha_len_03
// 
assign sha_len_03 = n0785;
// 
// sha_bytes_processed_03
// 
assign sha_bytes_processed_03 = n0918;
// 
// sha_wraddr_03
// 
assign sha_wraddr_03 = n0923;
// 
// dataout_03
// 
assign n0974 = 16'hfe0b;
assign n0975 = ( n0974 == addrin );
assign n0976 = ( n0975 && n0507 );
assign n0977 = ( n0976 ) ? ( sha_state ) : ( n0695 );
assign n0978 = ( n0672 ) ? ( n0977 ) : ( n0697 );
assign n0979 = ( n0502 ) ? ( n0943 ) : ( n0978 );
assign dataout_03 = n0979;
// 
// sha_rdaddr_03
// 
assign sha_rdaddr_03 = n0706;
// 
// aes_state_03
// 
assign n0980 = ( n0973 < aes_len );
assign n0981 = ( n0980 ) ? ( n0916 ) : ( n0661 );
assign n0982 = ( n0955 ) ? ( n0981 ) : ( n0964 );
assign aes_state_03 = n0982;
// 
// sha_state_03
// 
assign sha_state_03 = n0917;
// 
// sha_digest_03
// 
assign n0983 = { ( input_sha_func_11 ), ( input_sha_func_12 ), ( input_sha_func_13 ) };
assign n0984 = ( n0930 ) ? ( n0983 ) : ( sha_digest );
assign n0985 = ( n0928 ) ? ( n0984 ) : ( sha_digest );
assign n0986 = ( n0924 ) ? ( n0926 ) : ( n0985 );
assign sha_digest_03 = n0986;
assign n0987 = ( n0939 && n0930 );
assign n0988 = ( n0987 && n0955 );
assign n0989 = !( n0930 );
assign n0990 = ( n0939 && n0989 );
assign n0991 = ( n0990 && n0955 );
assign n0992 = !( n0938 );
assign n0993 = ( 1 && n0992 );
assign n0994 = ( n0993 && n0930 );
assign n0995 = ( n0994 && n0955 );
assign n0996 = ( n0993 && n0989 );
assign n0997 = ( n0996 && n0955 );
assign n0998 = ( nondet_memwrite_choice_103 ) ? ( n0997 ) : ( n0997 );
assign n0999 = ( nondet_memwrite_choice_102 ) ? ( n0997 ) : ( n0998 );
assign n1000 = ( nondet_memwrite_choice_101 ) ? ( n0997 ) : ( n0999 );
assign n1001 = ( nondet_memwrite_choice_100 ) ? ( n0997 ) : ( n1000 );
assign n1002 = ( nondet_memwrite_choice_99 ) ? ( n0997 ) : ( n1001 );
assign n1003 = ( nondet_memwrite_choice_98 ) ? ( n0997 ) : ( n1002 );
assign n1004 = ( nondet_memwrite_choice_97 ) ? ( n0997 ) : ( n1003 );
assign n1005 = ( nondet_memwrite_choice_96 ) ? ( n0997 ) : ( n1004 );
assign n1006 = ( nondet_memwrite_choice_95 ) ? ( n0997 ) : ( n1005 );
assign n1007 = ( nondet_memwrite_choice_94 ) ? ( n0997 ) : ( n1006 );
assign n1008 = ( nondet_memwrite_choice_93 ) ? ( n0997 ) : ( n1007 );
assign n1009 = ( nondet_memwrite_choice_92 ) ? ( n0997 ) : ( n1008 );
assign n1010 = ( nondet_memwrite_choice_91 ) ? ( n0997 ) : ( n1009 );
assign n1011 = ( nondet_memwrite_choice_90 ) ? ( n0997 ) : ( n1010 );
assign n1012 = ( nondet_memwrite_choice_89 ) ? ( n0997 ) : ( n1011 );
assign n1013 = ( nondet_memwrite_choice_88 ) ? ( n0995 ) : ( n1012 );
assign n1014 = ( nondet_memwrite_choice_87 ) ? ( n0995 ) : ( n1013 );
assign n1015 = ( nondet_memwrite_choice_86 ) ? ( n0995 ) : ( n1014 );
assign n1016 = ( nondet_memwrite_choice_85 ) ? ( n0995 ) : ( n1015 );
assign n1017 = ( nondet_memwrite_choice_84 ) ? ( n0995 ) : ( n1016 );
assign n1018 = ( nondet_memwrite_choice_83 ) ? ( n0995 ) : ( n1017 );
assign n1019 = ( nondet_memwrite_choice_82 ) ? ( n0995 ) : ( n1018 );
assign n1020 = ( nondet_memwrite_choice_81 ) ? ( n0995 ) : ( n1019 );
assign n1021 = ( nondet_memwrite_choice_80 ) ? ( n0995 ) : ( n1020 );
assign n1022 = ( nondet_memwrite_choice_79 ) ? ( n0995 ) : ( n1021 );
assign n1023 = ( nondet_memwrite_choice_78 ) ? ( n0995 ) : ( n1022 );
assign n1024 = ( nondet_memwrite_choice_77 ) ? ( n0995 ) : ( n1023 );
assign n1025 = ( nondet_memwrite_choice_76 ) ? ( n0995 ) : ( n1024 );
assign n1026 = ( nondet_memwrite_choice_75 ) ? ( n0995 ) : ( n1025 );
assign n1027 = ( nondet_memwrite_choice_74 ) ? ( n0995 ) : ( n1026 );
assign n1028 = ( nondet_memwrite_choice_73 ) ? ( n0995 ) : ( n1027 );
assign n1029 = ( nondet_memwrite_choice_72 ) ? ( n0994 ) : ( n1028 );
assign n1030 = ( nondet_memwrite_choice_71 ) ? ( n0994 ) : ( n1029 );
assign n1031 = ( nondet_memwrite_choice_70 ) ? ( n0994 ) : ( n1030 );
assign n1032 = ( nondet_memwrite_choice_69 ) ? ( n0994 ) : ( n1031 );
assign n1033 = ( nondet_memwrite_choice_68 ) ? ( n0994 ) : ( n1032 );
assign n1034 = ( nondet_memwrite_choice_67 ) ? ( n0994 ) : ( n1033 );
assign n1035 = ( nondet_memwrite_choice_66 ) ? ( n0994 ) : ( n1034 );
assign n1036 = ( nondet_memwrite_choice_65 ) ? ( n0994 ) : ( n1035 );
assign n1037 = ( nondet_memwrite_choice_64 ) ? ( n0994 ) : ( n1036 );
assign n1038 = ( nondet_memwrite_choice_63 ) ? ( n0994 ) : ( n1037 );
assign n1039 = ( nondet_memwrite_choice_62 ) ? ( n0994 ) : ( n1038 );
assign n1040 = ( nondet_memwrite_choice_61 ) ? ( n0994 ) : ( n1039 );
assign n1041 = ( nondet_memwrite_choice_60 ) ? ( n0994 ) : ( n1040 );
assign n1042 = ( nondet_memwrite_choice_59 ) ? ( n0994 ) : ( n1041 );
assign n1043 = ( nondet_memwrite_choice_58 ) ? ( n0994 ) : ( n1042 );
assign n1044 = ( nondet_memwrite_choice_57 ) ? ( n0994 ) : ( n1043 );
assign n1045 = ( nondet_memwrite_choice_56 ) ? ( n0994 ) : ( n1044 );
assign n1046 = ( nondet_memwrite_choice_55 ) ? ( n0994 ) : ( n1045 );
assign n1047 = ( nondet_memwrite_choice_54 ) ? ( n0994 ) : ( n1046 );
assign n1048 = ( nondet_memwrite_choice_53 ) ? ( n0994 ) : ( n1047 );
assign n1049 = ( nondet_memwrite_choice_52 ) ? ( n0991 ) : ( n1048 );
assign n1050 = ( nondet_memwrite_choice_51 ) ? ( n0991 ) : ( n1049 );
assign n1051 = ( nondet_memwrite_choice_50 ) ? ( n0991 ) : ( n1050 );
assign n1052 = ( nondet_memwrite_choice_49 ) ? ( n0991 ) : ( n1051 );
assign n1053 = ( nondet_memwrite_choice_48 ) ? ( n0991 ) : ( n1052 );
assign n1054 = ( nondet_memwrite_choice_47 ) ? ( n0991 ) : ( n1053 );
assign n1055 = ( nondet_memwrite_choice_46 ) ? ( n0991 ) : ( n1054 );
assign n1056 = ( nondet_memwrite_choice_45 ) ? ( n0991 ) : ( n1055 );
assign n1057 = ( nondet_memwrite_choice_44 ) ? ( n0991 ) : ( n1056 );
assign n1058 = ( nondet_memwrite_choice_43 ) ? ( n0991 ) : ( n1057 );
assign n1059 = ( nondet_memwrite_choice_42 ) ? ( n0991 ) : ( n1058 );
assign n1060 = ( nondet_memwrite_choice_41 ) ? ( n0991 ) : ( n1059 );
assign n1061 = ( nondet_memwrite_choice_40 ) ? ( n0991 ) : ( n1060 );
assign n1062 = ( nondet_memwrite_choice_39 ) ? ( n0991 ) : ( n1061 );
assign n1063 = ( nondet_memwrite_choice_38 ) ? ( n0991 ) : ( n1062 );
assign n1064 = ( nondet_memwrite_choice_37 ) ? ( n0991 ) : ( n1063 );
assign n1065 = ( nondet_memwrite_choice_36 ) ? ( n0988 ) : ( n1064 );
assign n1066 = ( nondet_memwrite_choice_35 ) ? ( n0988 ) : ( n1065 );
assign n1067 = ( nondet_memwrite_choice_34 ) ? ( n0988 ) : ( n1066 );
assign n1068 = ( nondet_memwrite_choice_33 ) ? ( n0988 ) : ( n1067 );
assign n1069 = ( nondet_memwrite_choice_32 ) ? ( n0988 ) : ( n1068 );
assign n1070 = ( nondet_memwrite_choice_31 ) ? ( n0988 ) : ( n1069 );
assign n1071 = ( nondet_memwrite_choice_30 ) ? ( n0988 ) : ( n1070 );
assign n1072 = ( nondet_memwrite_choice_29 ) ? ( n0988 ) : ( n1071 );
assign n1073 = ( nondet_memwrite_choice_28 ) ? ( n0988 ) : ( n1072 );
assign n1074 = ( nondet_memwrite_choice_27 ) ? ( n0988 ) : ( n1073 );
assign n1075 = ( nondet_memwrite_choice_26 ) ? ( n0988 ) : ( n1074 );
assign n1076 = ( nondet_memwrite_choice_25 ) ? ( n0988 ) : ( n1075 );
assign n1077 = ( nondet_memwrite_choice_24 ) ? ( n0988 ) : ( n1076 );
assign n1078 = ( nondet_memwrite_choice_23 ) ? ( n0988 ) : ( n1077 );
assign n1079 = ( nondet_memwrite_choice_22 ) ? ( n0988 ) : ( n1078 );
assign n1080 = ( nondet_memwrite_choice_21 ) ? ( n0988 ) : ( n1079 );
assign n1081 = ( nondet_memwrite_choice_20 ) ? ( n0987 ) : ( n1080 );
assign n1082 = ( nondet_memwrite_choice_19 ) ? ( n0987 ) : ( n1081 );
assign n1083 = ( nondet_memwrite_choice_18 ) ? ( n0987 ) : ( n1082 );
assign n1084 = ( nondet_memwrite_choice_17 ) ? ( n0987 ) : ( n1083 );
assign n1085 = ( nondet_memwrite_choice_16 ) ? ( n0987 ) : ( n1084 );
assign n1086 = ( nondet_memwrite_choice_15 ) ? ( n0987 ) : ( n1085 );
assign n1087 = ( nondet_memwrite_choice_14 ) ? ( n0987 ) : ( n1086 );
assign n1088 = ( nondet_memwrite_choice_13 ) ? ( n0987 ) : ( n1087 );
assign n1089 = ( nondet_memwrite_choice_12 ) ? ( n0987 ) : ( n1088 );
assign n1090 = ( nondet_memwrite_choice_11 ) ? ( n0987 ) : ( n1089 );
assign n1091 = ( nondet_memwrite_choice_10 ) ? ( n0987 ) : ( n1090 );
assign n1092 = ( nondet_memwrite_choice_9 ) ? ( n0987 ) : ( n1091 );
assign n1093 = ( nondet_memwrite_choice_8 ) ? ( n0987 ) : ( n1092 );
assign n1094 = ( nondet_memwrite_choice_7 ) ? ( n0987 ) : ( n1093 );
assign n1095 = ( nondet_memwrite_choice_6 ) ? ( n0987 ) : ( n1094 );
assign n1096 = ( nondet_memwrite_choice_5 ) ? ( n0987 ) : ( n1095 );
assign n1097 = ( nondet_memwrite_choice_4 ) ? ( n0987 ) : ( n1096 );
assign n1098 = ( nondet_memwrite_choice_3 ) ? ( n0987 ) : ( n1097 );
assign n1099 = ( nondet_memwrite_choice_2 ) ? ( n0987 ) : ( n1098 );
assign n1100 = ( nondet_memwrite_choice_1 ) ? ( n0987 ) : ( n1099 );
assign n1101 = ( nondet_memwrite_choice_0 ) ? ( n0939 ) : ( n1100 );
assign WR_XRAM_EN_03 = n1101;
assign n1102 = ( sha_wraddr + n0395 );
assign n1103 = ( sha_wraddr + n0401 );
assign n1104 = ( sha_wraddr + n0407 );
assign n1105 = ( sha_wraddr + n0413 );
assign n1106 = ( sha_wraddr + n0418 );
assign n1107 = ( sha_wraddr + n0423 );
assign n1108 = ( sha_wraddr + n0428 );
assign n1109 = ( sha_wraddr + n0433 );
assign n1110 = ( sha_wraddr + n0438 );
assign n1111 = ( sha_wraddr + n0443 );
assign n1112 = ( sha_wraddr + n0448 );
assign n1113 = ( sha_wraddr + n0453 );
assign n1114 = ( sha_wraddr + n0458 );
assign n1115 = ( sha_wraddr + n0463 );
assign n1116 = ( sha_wraddr + n0468 );
assign n1117 = ( sha_wraddr + n0473 );
assign n1118 = ( sha_wraddr + n0478 );
assign n1119 = ( sha_wraddr + n0483 );
assign n1120 = ( sha_wraddr + n0488 );
assign n1121 = ( sha_wraddr + n0493 );
assign n1122 = ( nondet_memwrite_choice_103 ) ? ( n0199 ) : ( n0210 );
assign n1123 = ( nondet_memwrite_choice_102 ) ? ( n0188 ) : ( n1122 );
assign n1124 = ( nondet_memwrite_choice_101 ) ? ( n0177 ) : ( n1123 );
assign n1125 = ( nondet_memwrite_choice_100 ) ? ( n0166 ) : ( n1124 );
assign n1126 = ( nondet_memwrite_choice_99 ) ? ( n0155 ) : ( n1125 );
assign n1127 = ( nondet_memwrite_choice_98 ) ? ( n0144 ) : ( n1126 );
assign n1128 = ( nondet_memwrite_choice_97 ) ? ( n0133 ) : ( n1127 );
assign n1129 = ( nondet_memwrite_choice_96 ) ? ( n0122 ) : ( n1128 );
assign n1130 = ( nondet_memwrite_choice_95 ) ? ( n0111 ) : ( n1129 );
assign n1131 = ( nondet_memwrite_choice_94 ) ? ( n0100 ) : ( n1130 );
assign n1132 = ( nondet_memwrite_choice_93 ) ? ( n0089 ) : ( n1131 );
assign n1133 = ( nondet_memwrite_choice_92 ) ? ( n0078 ) : ( n1132 );
assign n1134 = ( nondet_memwrite_choice_91 ) ? ( n0067 ) : ( n1133 );
assign n1135 = ( nondet_memwrite_choice_90 ) ? ( n0056 ) : ( n1134 );
assign n1136 = ( nondet_memwrite_choice_89 ) ? ( n0034 ) : ( n1135 );
assign n1137 = ( nondet_memwrite_choice_88 ) ? ( n0210 ) : ( n1136 );
assign n1138 = ( nondet_memwrite_choice_87 ) ? ( n0199 ) : ( n1137 );
assign n1139 = ( nondet_memwrite_choice_86 ) ? ( n0188 ) : ( n1138 );
assign n1140 = ( nondet_memwrite_choice_85 ) ? ( n0177 ) : ( n1139 );
assign n1141 = ( nondet_memwrite_choice_84 ) ? ( n0166 ) : ( n1140 );
assign n1142 = ( nondet_memwrite_choice_83 ) ? ( n0155 ) : ( n1141 );
assign n1143 = ( nondet_memwrite_choice_82 ) ? ( n0144 ) : ( n1142 );
assign n1144 = ( nondet_memwrite_choice_81 ) ? ( n0133 ) : ( n1143 );
assign n1145 = ( nondet_memwrite_choice_80 ) ? ( n0122 ) : ( n1144 );
assign n1146 = ( nondet_memwrite_choice_79 ) ? ( n0111 ) : ( n1145 );
assign n1147 = ( nondet_memwrite_choice_78 ) ? ( n0100 ) : ( n1146 );
assign n1148 = ( nondet_memwrite_choice_77 ) ? ( n0089 ) : ( n1147 );
assign n1149 = ( nondet_memwrite_choice_76 ) ? ( n0078 ) : ( n1148 );
assign n1150 = ( nondet_memwrite_choice_75 ) ? ( n0067 ) : ( n1149 );
assign n1151 = ( nondet_memwrite_choice_74 ) ? ( n0056 ) : ( n1150 );
assign n1152 = ( nondet_memwrite_choice_73 ) ? ( n0034 ) : ( n1151 );
assign n1153 = ( nondet_memwrite_choice_72 ) ? ( n1121 ) : ( n1152 );
assign n1154 = ( nondet_memwrite_choice_71 ) ? ( n1120 ) : ( n1153 );
assign n1155 = ( nondet_memwrite_choice_70 ) ? ( n1119 ) : ( n1154 );
assign n1156 = ( nondet_memwrite_choice_69 ) ? ( n1118 ) : ( n1155 );
assign n1157 = ( nondet_memwrite_choice_68 ) ? ( n1117 ) : ( n1156 );
assign n1158 = ( nondet_memwrite_choice_67 ) ? ( n1116 ) : ( n1157 );
assign n1159 = ( nondet_memwrite_choice_66 ) ? ( n1115 ) : ( n1158 );
assign n1160 = ( nondet_memwrite_choice_65 ) ? ( n1114 ) : ( n1159 );
assign n1161 = ( nondet_memwrite_choice_64 ) ? ( n1113 ) : ( n1160 );
assign n1162 = ( nondet_memwrite_choice_63 ) ? ( n1112 ) : ( n1161 );
assign n1163 = ( nondet_memwrite_choice_62 ) ? ( n1111 ) : ( n1162 );
assign n1164 = ( nondet_memwrite_choice_61 ) ? ( n1110 ) : ( n1163 );
assign n1165 = ( nondet_memwrite_choice_60 ) ? ( n1109 ) : ( n1164 );
assign n1166 = ( nondet_memwrite_choice_59 ) ? ( n1108 ) : ( n1165 );
assign n1167 = ( nondet_memwrite_choice_58 ) ? ( n1107 ) : ( n1166 );
assign n1168 = ( nondet_memwrite_choice_57 ) ? ( n1106 ) : ( n1167 );
assign n1169 = ( nondet_memwrite_choice_56 ) ? ( n1105 ) : ( n1168 );
assign n1170 = ( nondet_memwrite_choice_55 ) ? ( n1104 ) : ( n1169 );
assign n1171 = ( nondet_memwrite_choice_54 ) ? ( n1103 ) : ( n1170 );
assign n1172 = ( nondet_memwrite_choice_53 ) ? ( n1102 ) : ( n1171 );
assign n1173 = ( nondet_memwrite_choice_52 ) ? ( n0210 ) : ( n1172 );
assign n1174 = ( nondet_memwrite_choice_51 ) ? ( n0199 ) : ( n1173 );
assign n1175 = ( nondet_memwrite_choice_50 ) ? ( n0188 ) : ( n1174 );
assign n1176 = ( nondet_memwrite_choice_49 ) ? ( n0177 ) : ( n1175 );
assign n1177 = ( nondet_memwrite_choice_48 ) ? ( n0166 ) : ( n1176 );
assign n1178 = ( nondet_memwrite_choice_47 ) ? ( n0155 ) : ( n1177 );
assign n1179 = ( nondet_memwrite_choice_46 ) ? ( n0144 ) : ( n1178 );
assign n1180 = ( nondet_memwrite_choice_45 ) ? ( n0133 ) : ( n1179 );
assign n1181 = ( nondet_memwrite_choice_44 ) ? ( n0122 ) : ( n1180 );
assign n1182 = ( nondet_memwrite_choice_43 ) ? ( n0111 ) : ( n1181 );
assign n1183 = ( nondet_memwrite_choice_42 ) ? ( n0100 ) : ( n1182 );
assign n1184 = ( nondet_memwrite_choice_41 ) ? ( n0089 ) : ( n1183 );
assign n1185 = ( nondet_memwrite_choice_40 ) ? ( n0078 ) : ( n1184 );
assign n1186 = ( nondet_memwrite_choice_39 ) ? ( n0067 ) : ( n1185 );
assign n1187 = ( nondet_memwrite_choice_38 ) ? ( n0056 ) : ( n1186 );
assign n1188 = ( nondet_memwrite_choice_37 ) ? ( n0034 ) : ( n1187 );
assign n1189 = ( nondet_memwrite_choice_36 ) ? ( n0210 ) : ( n1188 );
assign n1190 = ( nondet_memwrite_choice_35 ) ? ( n0199 ) : ( n1189 );
assign n1191 = ( nondet_memwrite_choice_34 ) ? ( n0188 ) : ( n1190 );
assign n1192 = ( nondet_memwrite_choice_33 ) ? ( n0177 ) : ( n1191 );
assign n1193 = ( nondet_memwrite_choice_32 ) ? ( n0166 ) : ( n1192 );
assign n1194 = ( nondet_memwrite_choice_31 ) ? ( n0155 ) : ( n1193 );
assign n1195 = ( nondet_memwrite_choice_30 ) ? ( n0144 ) : ( n1194 );
assign n1196 = ( nondet_memwrite_choice_29 ) ? ( n0133 ) : ( n1195 );
assign n1197 = ( nondet_memwrite_choice_28 ) ? ( n0122 ) : ( n1196 );
assign n1198 = ( nondet_memwrite_choice_27 ) ? ( n0111 ) : ( n1197 );
assign n1199 = ( nondet_memwrite_choice_26 ) ? ( n0100 ) : ( n1198 );
assign n1200 = ( nondet_memwrite_choice_25 ) ? ( n0089 ) : ( n1199 );
assign n1201 = ( nondet_memwrite_choice_24 ) ? ( n0078 ) : ( n1200 );
assign n1202 = ( nondet_memwrite_choice_23 ) ? ( n0067 ) : ( n1201 );
assign n1203 = ( nondet_memwrite_choice_22 ) ? ( n0056 ) : ( n1202 );
assign n1204 = ( nondet_memwrite_choice_21 ) ? ( n0034 ) : ( n1203 );
assign n1205 = ( nondet_memwrite_choice_20 ) ? ( n1121 ) : ( n1204 );
assign n1206 = ( nondet_memwrite_choice_19 ) ? ( n1120 ) : ( n1205 );
assign n1207 = ( nondet_memwrite_choice_18 ) ? ( n1119 ) : ( n1206 );
assign n1208 = ( nondet_memwrite_choice_17 ) ? ( n1118 ) : ( n1207 );
assign n1209 = ( nondet_memwrite_choice_16 ) ? ( n1117 ) : ( n1208 );
assign n1210 = ( nondet_memwrite_choice_15 ) ? ( n1116 ) : ( n1209 );
assign n1211 = ( nondet_memwrite_choice_14 ) ? ( n1115 ) : ( n1210 );
assign n1212 = ( nondet_memwrite_choice_13 ) ? ( n1114 ) : ( n1211 );
assign n1213 = ( nondet_memwrite_choice_12 ) ? ( n1113 ) : ( n1212 );
assign n1214 = ( nondet_memwrite_choice_11 ) ? ( n1112 ) : ( n1213 );
assign n1215 = ( nondet_memwrite_choice_10 ) ? ( n1111 ) : ( n1214 );
assign n1216 = ( nondet_memwrite_choice_9 ) ? ( n1110 ) : ( n1215 );
assign n1217 = ( nondet_memwrite_choice_8 ) ? ( n1109 ) : ( n1216 );
assign n1218 = ( nondet_memwrite_choice_7 ) ? ( n1108 ) : ( n1217 );
assign n1219 = ( nondet_memwrite_choice_6 ) ? ( n1107 ) : ( n1218 );
assign n1220 = ( nondet_memwrite_choice_5 ) ? ( n1106 ) : ( n1219 );
assign n1221 = ( nondet_memwrite_choice_4 ) ? ( n1105 ) : ( n1220 );
assign n1222 = ( nondet_memwrite_choice_3 ) ? ( n1104 ) : ( n1221 );
assign n1223 = ( nondet_memwrite_choice_2 ) ? ( n1103 ) : ( n1222 );
assign n1224 = ( nondet_memwrite_choice_1 ) ? ( n1102 ) : ( n1223 );
assign n1225 = ( nondet_memwrite_choice_0 ) ? ( addrin ) : ( n1224 );
assign WR_XRAM_ADDR_03 = n1225;
// 
// dataout_04
// 
assign n1226 = 16'hff08;
assign n1227 = ( n1226 == addrin );
assign n1228 = ( n1227 && n0507 );
assign n1229 = ( n1228 ) ? ( aes_state ) : ( n0666 );
assign n1230 = 16'hfe01;
assign n1231 = ( n1230 == addrin );
assign n1232 = ( n1231 && n0507 );
assign n1233 = ( n1232 ) ? ( sha_state ) : ( n0695 );
assign n1234 = ( n0672 ) ? ( n1233 ) : ( n0697 );
assign n1235 = ( n0502 ) ? ( n1229 ) : ( n1234 );
assign dataout_04 = n1235;
// 
// aes_addr_04
// 
assign aes_addr_04 = n0713;
// 
// aes_ctr_04
// 
assign aes_ctr_04 = n0774;
// 
// aes_bytes_processed_04
// 
assign aes_bytes_processed_04 = n0780;
// 
// aes_key1_04
// 
assign aes_key1_04 = n0846;
// 
// aes_key0_04
// 
assign aes_key0_04 = n0907;
// 
// aes_len_04
// 
assign aes_len_04 = n0912;
// 
// sha_bytes_processed_04
// 
assign sha_bytes_processed_04 = n0918;
// 
// sha_digest_04
// 
assign n1236 = { ( input_sha_func_14 ), ( input_sha_func_15 ), ( input_sha_func_16 ) };
assign n1237 = ( n0930 ) ? ( n1236 ) : ( sha_digest );
assign n1238 = ( n0928 ) ? ( n1237 ) : ( sha_digest );
assign n1239 = ( n0924 ) ? ( n0926 ) : ( n1238 );
assign sha_digest_04 = n1239;
// 
// sha_read_data_04
// 
assign n1240 = { ( RD_xram_1 ), ( RD_xram_2 ), ( RD_xram_3 ), ( RD_xram_4 ), ( RD_xram_5 ), ( RD_xram_6 ), ( RD_xram_7 ), ( RD_xram_8 ), ( RD_xram_9 ), ( RD_xram_10 ), ( RD_xram_11 ), ( RD_xram_12 ), ( RD_xram_13 ), ( RD_xram_14 ), ( RD_xram_15 ), ( RD_xram_16 ), ( RD_xram_17 ), ( RD_xram_18 ), ( RD_xram_19 ), ( RD_xram_20 ), ( RD_xram_21 ), ( RD_xram_22 ), ( RD_xram_23 ), ( RD_xram_24 ), ( RD_xram_25 ), ( RD_xram_26 ), ( RD_xram_27 ), ( RD_xram_28 ), ( RD_xram_29 ), ( RD_xram_30 ), ( RD_xram_31 ), ( RD_xram_32 ), ( RD_xram_33 ), ( RD_xram_34 ), ( RD_xram_35 ), ( RD_xram_36 ), ( RD_xram_37 ), ( RD_xram_38 ), ( RD_xram_39 ), ( RD_xram_40 ), ( RD_xram_41 ), ( RD_xram_42 ), ( RD_xram_43 ), ( RD_xram_44 ), ( RD_xram_45 ), ( RD_xram_46 ), ( RD_xram_47 ), ( RD_xram_48 ), ( RD_xram_49 ), ( RD_xram_50 ), ( RD_xram_51 ), ( RD_xram_52 ), ( RD_xram_53 ), ( RD_xram_54 ), ( RD_xram_55 ), ( RD_xram_56 ), ( RD_xram_57 ), ( RD_xram_58 ), ( RD_xram_59 ), ( RD_xram_60 ), ( RD_xram_61 ), ( RD_xram_62 ), ( RD_xram_63 ), ( RD_xram_64 ) };
assign n1241 = ( n0930 ) ? ( n1240 ) : ( sha_read_data );
assign sha_read_data_04 = n1241;
// 
// xram_04
// 
// 
// aes_state_04
// 
assign aes_state_04 = n0935;
// 
// sha_state_04
// 
assign n1242 = ( n0930 ) ? ( n0927 ) : ( n0916 );
assign sha_state_04 = n1242;
assign WR_XRAM_EN_04 = n0939;
assign WR_XRAM_ADDR_04 = addrin;
// 
// xram_05
// 
// 
// dataout_05
// 
assign n1243 = ( n0502 ) ? ( n0943 ) : ( n1234 );
assign dataout_05 = n1243;
// 
// aes_bytes_processed_05
// 
assign aes_bytes_processed_05 = n0953;
// 
// aes_read_data_05
// 
assign aes_read_data_05 = n0957;
// 
// sha_bytes_processed_05
// 
assign sha_bytes_processed_05 = n0918;
// 
// sha_digest_05
// 
assign n1244 = { ( input_sha_func_17 ), ( input_sha_func_18 ), ( input_sha_func_19 ) };
assign n1245 = ( n0930 ) ? ( n1244 ) : ( sha_digest );
assign n1246 = ( n0928 ) ? ( n1245 ) : ( sha_digest );
assign n1247 = ( n0924 ) ? ( n0926 ) : ( n1246 );
assign sha_digest_05 = n1247;
// 
// sha_read_data_05
// 
assign n1248 = { ( RD_xram_17 ), ( RD_xram_18 ), ( RD_xram_19 ), ( RD_xram_20 ), ( RD_xram_21 ), ( RD_xram_22 ), ( RD_xram_23 ), ( RD_xram_24 ), ( RD_xram_25 ), ( RD_xram_26 ), ( RD_xram_27 ), ( RD_xram_28 ), ( RD_xram_29 ), ( RD_xram_30 ), ( RD_xram_31 ), ( RD_xram_32 ), ( RD_xram_33 ), ( RD_xram_34 ), ( RD_xram_35 ), ( RD_xram_36 ), ( RD_xram_37 ), ( RD_xram_38 ), ( RD_xram_39 ), ( RD_xram_40 ), ( RD_xram_41 ), ( RD_xram_42 ), ( RD_xram_43 ), ( RD_xram_44 ), ( RD_xram_45 ), ( RD_xram_46 ), ( RD_xram_47 ), ( RD_xram_48 ), ( RD_xram_49 ), ( RD_xram_50 ), ( RD_xram_51 ), ( RD_xram_52 ), ( RD_xram_53 ), ( RD_xram_54 ), ( RD_xram_55 ), ( RD_xram_56 ), ( RD_xram_57 ), ( RD_xram_58 ), ( RD_xram_59 ), ( RD_xram_60 ), ( RD_xram_61 ), ( RD_xram_62 ), ( RD_xram_63 ), ( RD_xram_64 ), ( RD_xram_65 ), ( RD_xram_66 ), ( RD_xram_67 ), ( RD_xram_68 ), ( RD_xram_69 ), ( RD_xram_70 ), ( RD_xram_71 ), ( RD_xram_72 ), ( RD_xram_73 ), ( RD_xram_74 ), ( RD_xram_75 ), ( RD_xram_76 ), ( RD_xram_77 ), ( RD_xram_78 ), ( RD_xram_79 ), ( RD_xram_80 ) };
assign n1249 = ( n0930 ) ? ( n1248 ) : ( sha_read_data );
assign sha_read_data_05 = n1249;
// 
// aes_state_05
// 
assign aes_state_05 = n0962;
// 
// sha_state_05
// 
assign sha_state_05 = n1242;
assign WR_XRAM_EN_05 = n0939;
assign WR_XRAM_ADDR_05 = addrin;
// 
// dataout_06
// 
assign dataout_06 = n1243;
// 
// aes_bytes_processed_06
// 
assign aes_bytes_processed_06 = n0953;
// 
// sha_state_06
// 
assign sha_state_06 = n1242;
// 
// sha_bytes_processed_06
// 
assign sha_bytes_processed_06 = n0918;
// 
// sha_digest_06
// 
assign n1250 = { ( input_sha_func_20 ), ( input_sha_func_21 ), ( input_sha_func_22 ) };
assign n1251 = ( n0930 ) ? ( n1250 ) : ( sha_digest );
assign n1252 = ( n0928 ) ? ( n1251 ) : ( sha_digest );
assign n1253 = ( n0924 ) ? ( n0926 ) : ( n1252 );
assign sha_digest_06 = n1253;
// 
// sha_read_data_06
// 
assign sha_read_data_06 = n1241;
// 
// xram_06
// 
// 
// aes_state_06
// 
assign aes_state_06 = n0965;
// 
// aes_enc_data_06
// 
assign n1254 = { ( input_aes_func_23 ), ( input_aes_func_24 ) };
assign n1255 = ( n0955 ) ? ( n1254 ) : ( aes_enc_data );
assign aes_enc_data_06 = n1255;
assign WR_XRAM_EN_06 = n0939;
assign WR_XRAM_ADDR_06 = addrin;
// 
// aes_bytes_processed_07
// 
assign aes_bytes_processed_07 = n0973;
// 
// sha_bytes_processed_07
// 
assign sha_bytes_processed_07 = n0918;
// 
// dataout_07
// 
assign dataout_07 = n1243;
// 
// sha_read_data_07
// 
assign sha_read_data_07 = n1241;
// 
// xram_07
// 
// 
// aes_state_07
// 
assign aes_state_07 = n0982;
// 
// sha_state_07
// 
assign sha_state_07 = n1242;
// 
// sha_digest_07
// 
assign n1256 = { ( input_sha_func_25 ), ( input_sha_func_26 ), ( input_sha_func_27 ) };
assign n1257 = ( n0930 ) ? ( n1256 ) : ( sha_digest );
assign n1258 = ( n0928 ) ? ( n1257 ) : ( sha_digest );
assign n1259 = ( n0924 ) ? ( n0926 ) : ( n1258 );
assign sha_digest_07 = n1259;
assign WR_XRAM_EN_07 = n1101;
assign WR_XRAM_ADDR_07 = n1225;
// 
// aes_key0_08
// 
assign aes_key0_08 = n0907;
// 
// xram_08
// 
// 
// aes_addr_08
// 
assign aes_addr_08 = n0713;
// 
// aes_ctr_08
// 
assign aes_ctr_08 = n0774;
// 
// aes_bytes_processed_08
// 
assign aes_bytes_processed_08 = n0780;
// 
// aes_key1_08
// 
assign aes_key1_08 = n0846;
// 
// dataout_08
// 
assign n1260 = ( n0502 ) ? ( n0667 ) : ( n1234 );
assign dataout_08 = n1260;
// 
// aes_len_08
// 
assign aes_len_08 = n0912;
// 
// sha_state_08
// 
assign n1261 = 16'h40;
assign n1262 = ( sha_bytes_processed + n1261 );
assign n1263 = ( n0930 ) ? ( n1262 ) : ( sha_bytes_processed );
assign n1264 = ( n1263 < sha_len );
assign n1265 = ( n1264 ) ? ( n0916 ) : ( n0964 );
assign n1266 = ( n0930 ) ? ( n1265 ) : ( n0927 );
assign sha_state_08 = n1266;
// 
// sha_bytes_processed_08
// 
assign sha_bytes_processed_08 = n1263;
// 
// sha_digest_08
// 
assign n1267 = { ( input_sha_func_28 ), ( input_sha_func_29 ), ( input_sha_func_30 ) };
assign n1268 = ( n0930 ) ? ( n1267 ) : ( sha_digest );
assign n1269 = ( n0928 ) ? ( n1268 ) : ( sha_digest );
assign n1270 = ( n0924 ) ? ( n0926 ) : ( n1269 );
assign sha_digest_08 = n1270;
// 
// aes_state_08
// 
assign aes_state_08 = n0935;
assign WR_XRAM_EN_08 = n0939;
assign WR_XRAM_ADDR_08 = addrin;
// 
// dataout_09
// 
assign dataout_09 = n1243;
// 
// xram_09
// 
// 
// aes_bytes_processed_09
// 
assign aes_bytes_processed_09 = n0953;
// 
// aes_read_data_09
// 
assign aes_read_data_09 = n0957;
// 
// sha_state_09
// 
assign sha_state_09 = n1266;
// 
// sha_bytes_processed_09
// 
assign sha_bytes_processed_09 = n1263;
// 
// sha_digest_09
// 
assign n1271 = { ( input_sha_func_31 ), ( input_sha_func_32 ), ( input_sha_func_33 ) };
assign n1272 = ( n0930 ) ? ( n1271 ) : ( sha_digest );
assign n1273 = ( n0928 ) ? ( n1272 ) : ( sha_digest );
assign n1274 = ( n0924 ) ? ( n0926 ) : ( n1273 );
assign sha_digest_09 = n1274;
// 
// aes_state_09
// 
assign aes_state_09 = n0962;
assign WR_XRAM_EN_09 = n0939;
assign WR_XRAM_ADDR_09 = addrin;
// 
// sha_digest_0a
// 
assign n1275 = { ( input_sha_func_34 ), ( input_sha_func_35 ), ( input_sha_func_36 ) };
assign n1276 = ( n0930 ) ? ( n1275 ) : ( sha_digest );
assign n1277 = ( n0928 ) ? ( n1276 ) : ( sha_digest );
assign n1278 = ( n0924 ) ? ( n0926 ) : ( n1277 );
assign sha_digest_0a = n1278;
// 
// aes_bytes_processed_0a
// 
assign aes_bytes_processed_0a = n0953;
// 
// sha_bytes_processed_0a
// 
assign sha_bytes_processed_0a = n1263;
// 
// dataout_0a
// 
assign dataout_0a = n1243;
// 
// xram_0a
// 
// 
// aes_state_0a
// 
assign aes_state_0a = n0965;
// 
// sha_state_0a
// 
assign sha_state_0a = n1266;
// 
// aes_enc_data_0a
// 
assign n1279 = { ( input_aes_func_37 ), ( input_aes_func_38 ) };
assign n1280 = ( n0955 ) ? ( n1279 ) : ( aes_enc_data );
assign aes_enc_data_0a = n1280;
assign WR_XRAM_EN_0a = n0939;
assign WR_XRAM_ADDR_0a = addrin;
// 
// sha_digest_0b
// 
assign n1281 = { ( input_sha_func_39 ), ( input_sha_func_40 ), ( input_sha_func_41 ) };
assign n1282 = ( n0930 ) ? ( n1281 ) : ( sha_digest );
assign n1283 = ( n0928 ) ? ( n1282 ) : ( sha_digest );
assign n1284 = ( n0924 ) ? ( n0926 ) : ( n1283 );
assign sha_digest_0b = n1284;
// 
// xram_0b
// 
// 
// aes_bytes_processed_0b
// 
assign aes_bytes_processed_0b = n0973;
// 
// sha_state_0b
// 
assign sha_state_0b = n1266;
// 
// sha_bytes_processed_0b
// 
assign sha_bytes_processed_0b = n1263;
// 
// dataout_0b
// 
assign dataout_0b = n1243;
// 
// aes_state_0b
// 
assign aes_state_0b = n0982;
assign WR_XRAM_EN_0b = n1101;
assign WR_XRAM_ADDR_0b = n1225;
// 
// aes_key0_0c
// 
assign aes_key0_0c = n0907;
// 
// xram_0c
// 
// 
// aes_addr_0c
// 
assign aes_addr_0c = n0713;
// 
// aes_key1_0c
// 
assign aes_key1_0c = n0846;
// 
// aes_bytes_processed_0c
// 
assign aes_bytes_processed_0c = n0780;
// 
// dataout_0c
// 
assign dataout_0c = n1243;
// 
// aes_len_0c
// 
assign aes_len_0c = n0912;
// 
// sha_bytes_processed_0c
// 
assign sha_bytes_processed_0c = n0918;
// 
// sha_digest_0c
// 
assign n1285 = { ( input_sha_func_42 ), ( input_sha_func_43 ), ( input_sha_func_44 ) };
assign n1286 = ( n0930 ) ? ( n1285 ) : ( sha_digest );
assign n1287 = ( n0928 ) ? ( n1286 ) : ( sha_digest );
assign n1288 = ( n0924 ) ? ( n0926 ) : ( n1287 );
assign sha_digest_0c = n1288;
// 
// aes_ctr_0c
// 
assign aes_ctr_0c = n0774;
// 
// aes_state_0c
// 
assign aes_state_0c = n0935;
// 
// sha_state_0c
// 
assign n1289 = ( n0930 ) ? ( n0661 ) : ( n0964 );
assign sha_state_0c = n1289;
assign WR_XRAM_EN_0c = n0939;
assign WR_XRAM_ADDR_0c = addrin;
// 
// xram_0d
// 
// 
// aes_bytes_processed_0d
// 
assign aes_bytes_processed_0d = n0953;
// 
// aes_read_data_0d
// 
assign n1290 = { ( RD_xram_0 ), ( RD_xram_1 ), ( RD_xram_2 ), ( RD_xram_3 ), ( RD_xram_4 ), ( RD_xram_5 ), ( RD_xram_6 ), ( RD_xram_7 ), ( RD_xram_8 ), ( RD_xram_9 ), ( RD_xram_10 ), ( RD_xram_11 ), ( RD_xram_12 ), ( RD_xram_13 ), ( RD_xram_14 ), ( RD_xram_15 ) };
assign n1291 = ( n0955 ) ? ( n1290 ) : ( aes_read_data );
assign aes_read_data_0d = n1291;
// 
// dataout_0d
// 
assign n1292 = ( n0507 ) ? ( RD_xram_16 ) : ( n0661 );
assign n1293 = ( n0672 ) ? ( n1233 ) : ( n1292 );
assign n1294 = ( n0502 ) ? ( n0943 ) : ( n1293 );
assign dataout_0d = n1294;
// 
// sha_state_0d
// 
assign sha_state_0d = n1289;
// 
// sha_bytes_processed_0d
// 
assign sha_bytes_processed_0d = n0918;
// 
// sha_digest_0d
// 
assign n1295 = { ( input_sha_func_45 ), ( input_sha_func_46 ), ( input_sha_func_47 ) };
assign n1296 = ( n0930 ) ? ( n1295 ) : ( sha_digest );
assign n1297 = ( n0928 ) ? ( n1296 ) : ( sha_digest );
assign n1298 = ( n0924 ) ? ( n0926 ) : ( n1297 );
assign sha_digest_0d = n1298;
// 
// aes_state_0d
// 
assign aes_state_0d = n0962;
assign WR_XRAM_EN_0d = n1101;
assign WR_XRAM_ADDR_0d = n1225;
// 
// aes_bytes_processed_0e
// 
assign aes_bytes_processed_0e = n0953;
// 
// dataout_0e
// 
assign dataout_0e = n1243;
// 
// sha_bytes_processed_0e
// 
assign sha_bytes_processed_0e = n0918;
// 
// sha_digest_0e
// 
assign n1299 = { ( input_sha_func_48 ), ( input_sha_func_49 ), ( input_sha_func_50 ) };
assign n1300 = ( n0930 ) ? ( n1299 ) : ( sha_digest );
assign n1301 = ( n0928 ) ? ( n1300 ) : ( sha_digest );
assign n1302 = ( n0924 ) ? ( n0926 ) : ( n1301 );
assign sha_digest_0e = n1302;
// 
// xram_0e
// 
// 
// aes_state_0e
// 
assign aes_state_0e = n0965;
// 
// sha_state_0e
// 
assign sha_state_0e = n1289;
// 
// aes_enc_data_0e
// 
assign n1303 = { ( input_aes_func_51 ), ( input_aes_func_52 ) };
assign n1304 = ( n0955 ) ? ( n1303 ) : ( aes_enc_data );
assign aes_enc_data_0e = n1304;
assign WR_XRAM_EN_0e = n0939;
assign WR_XRAM_ADDR_0e = addrin;
// 
// sha_digest_0f
// 
assign n1305 = { ( input_sha_func_53 ), ( input_sha_func_54 ), ( input_sha_func_55 ) };
assign n1306 = ( n0930 ) ? ( n1305 ) : ( sha_digest );
assign n1307 = ( n0928 ) ? ( n1306 ) : ( sha_digest );
assign n1308 = ( n0924 ) ? ( n0926 ) : ( n1307 );
assign sha_digest_0f = n1308;
// 
// xram_0f
// 
// 
// aes_bytes_processed_0f
// 
assign aes_bytes_processed_0f = n0973;
// 
// sha_bytes_processed_0f
// 
assign sha_bytes_processed_0f = n0918;
// 
// dataout_0f
// 
assign dataout_0f = n1243;
// 
// aes_state_0f
// 
assign aes_state_0f = n0982;
// 
// sha_state_0f
// 
assign sha_state_0f = n1289;
assign WR_XRAM_EN_0f = n1101;
assign WR_XRAM_ADDR_0f = n1225;
assign n1309 = ( n0003 == n0544 );
assign n1310 = ( n0003 == n0547 );
assign n1311 = ( n0003 == n0550 );
assign n1312 = ( n0003 == n0553 );
assign sha_read_data_next = 
  ( n1309 ) ? sha_read_data_04 : 
  ( n1310 ) ? sha_read_data_05 : 
  ( n1311 ) ? sha_read_data_06 : 
  ( n1312 ) ? sha_read_data_07 : 
  ( sha_read_data );
assign n1313 = ( n0003 == n0535 );
assign n1314 = ( n0003 == n0559 );
assign n1315 = ( n0003 == n0571 );
assign aes_read_data_next = 
  ( n1313 ) ? aes_read_data_01 : 
  ( n1310 ) ? aes_read_data_05 : 
  ( n1314 ) ? aes_read_data_09 : 
  ( n1315 ) ? aes_read_data_0d : 
  ( aes_read_data );
assign n1316 = ( n0003 == n0528 );
assign n1317 = ( n0003 == n0538 );
assign n1318 = ( n0003 == n0541 );
assign sha_rdaddr_next = 
  ( n1316 ) ? sha_rdaddr_00 : 
  ( n1313 ) ? sha_rdaddr_01 : 
  ( n1317 ) ? sha_rdaddr_02 : 
  ( n1318 ) ? sha_rdaddr_03 : 
  ( sha_rdaddr );
assign n1319 = ( n0003 == n0556 );
assign n1320 = ( n0003 == n0568 );
assign aes_addr_next = 
  ( n1316 ) ? aes_addr_00 : 
  ( n1309 ) ? aes_addr_04 : 
  ( n1319 ) ? aes_addr_08 : 
  ( n1320 ) ? aes_addr_0c : 
  ( aes_addr );
assign aes_ctr_next = 
  ( n1316 ) ? aes_ctr_00 : 
  ( n1309 ) ? aes_ctr_04 : 
  ( n1319 ) ? aes_ctr_08 : 
  ( n1320 ) ? aes_ctr_0c : 
  ( aes_ctr );
assign n1321 = ( n0003 == n0562 );
assign n1322 = ( n0003 == n0565 );
assign n1323 = ( n0003 == n0574 );
assign n1324 = 4'hf;
assign n1325 = ( n0003 == n1324 );
assign aes_bytes_processed_next = 
  ( n1316 ) ? aes_bytes_processed_00 : 
  ( n1313 ) ? aes_bytes_processed_01 : 
  ( n1317 ) ? aes_bytes_processed_02 : 
  ( n1318 ) ? aes_bytes_processed_03 : 
  ( n1309 ) ? aes_bytes_processed_04 : 
  ( n1310 ) ? aes_bytes_processed_05 : 
  ( n1311 ) ? aes_bytes_processed_06 : 
  ( n1312 ) ? aes_bytes_processed_07 : 
  ( n1319 ) ? aes_bytes_processed_08 : 
  ( n1314 ) ? aes_bytes_processed_09 : 
  ( n1321 ) ? aes_bytes_processed_0a : 
  ( n1322 ) ? aes_bytes_processed_0b : 
  ( n1320 ) ? aes_bytes_processed_0c : 
  ( n1315 ) ? aes_bytes_processed_0d : 
  ( n1323 ) ? aes_bytes_processed_0e : 
  ( n1325 ) ? aes_bytes_processed_0f : 
  ( aes_bytes_processed );
assign sha_len_next = 
  ( n1316 ) ? sha_len_00 : 
  ( n1313 ) ? sha_len_01 : 
  ( n1317 ) ? sha_len_02 : 
  ( n1318 ) ? sha_len_03 : 
  ( sha_len );
assign aes_key1_next = 
  ( n1316 ) ? aes_key1_00 : 
  ( n1309 ) ? aes_key1_04 : 
  ( n1319 ) ? aes_key1_08 : 
  ( n1320 ) ? aes_key1_0c : 
  ( aes_key1 );
assign aes_key0_next = 
  ( n1316 ) ? aes_key0_00 : 
  ( n1309 ) ? aes_key0_04 : 
  ( n1319 ) ? aes_key0_08 : 
  ( n1320 ) ? aes_key0_0c : 
  ( aes_key0 );
assign aes_len_next = 
  ( n1316 ) ? aes_len_00 : 
  ( n1309 ) ? aes_len_04 : 
  ( n1319 ) ? aes_len_08 : 
  ( n1320 ) ? aes_len_0c : 
  ( aes_len );
assign sha_bytes_processed_next = 
  ( n1316 ) ? sha_bytes_processed_00 : 
  ( n1313 ) ? sha_bytes_processed_01 : 
  ( n1317 ) ? sha_bytes_processed_02 : 
  ( n1318 ) ? sha_bytes_processed_03 : 
  ( n1309 ) ? sha_bytes_processed_04 : 
  ( n1310 ) ? sha_bytes_processed_05 : 
  ( n1311 ) ? sha_bytes_processed_06 : 
  ( n1312 ) ? sha_bytes_processed_07 : 
  ( n1319 ) ? sha_bytes_processed_08 : 
  ( n1314 ) ? sha_bytes_processed_09 : 
  ( n1321 ) ? sha_bytes_processed_0a : 
  ( n1322 ) ? sha_bytes_processed_0b : 
  ( n1320 ) ? sha_bytes_processed_0c : 
  ( n1315 ) ? sha_bytes_processed_0d : 
  ( n1323 ) ? sha_bytes_processed_0e : 
  ( n1325 ) ? sha_bytes_processed_0f : 
  ( sha_bytes_processed );
assign sha_wraddr_next = 
  ( n1316 ) ? sha_wraddr_00 : 
  ( n1313 ) ? sha_wraddr_01 : 
  ( n1317 ) ? sha_wraddr_02 : 
  ( n1318 ) ? sha_wraddr_03 : 
  ( sha_wraddr );
assign dataout_next = 
  ( n1316 ) ? dataout_00 : 
  ( n1313 ) ? dataout_01 : 
  ( n1317 ) ? dataout_02 : 
  ( n1318 ) ? dataout_03 : 
  ( n1309 ) ? dataout_04 : 
  ( n1310 ) ? dataout_05 : 
  ( n1311 ) ? dataout_06 : 
  ( n1312 ) ? dataout_07 : 
  ( n1319 ) ? dataout_08 : 
  ( n1314 ) ? dataout_09 : 
  ( n1321 ) ? dataout_0a : 
  ( n1322 ) ? dataout_0b : 
  ( n1320 ) ? dataout_0c : 
  ( n1315 ) ? dataout_0d : 
  ( n1323 ) ? dataout_0e : 
  ( n1325 ) ? dataout_0f : 
  ( dataout );
assign WR_XRAM_ADDR_next = 
  ( n1316 ) ? WR_XRAM_ADDR_00 : 
  ( n1313 ) ? WR_XRAM_ADDR_01 : 
  ( n1317 ) ? WR_XRAM_ADDR_02 : 
  ( n1318 ) ? WR_XRAM_ADDR_03 : 
  ( n1309 ) ? WR_XRAM_ADDR_04 : 
  ( n1310 ) ? WR_XRAM_ADDR_05 : 
  ( n1311 ) ? WR_XRAM_ADDR_06 : 
  ( n1312 ) ? WR_XRAM_ADDR_07 : 
  ( n1319 ) ? WR_XRAM_ADDR_08 : 
  ( n1314 ) ? WR_XRAM_ADDR_09 : 
  ( n1321 ) ? WR_XRAM_ADDR_0a : 
  ( n1322 ) ? WR_XRAM_ADDR_0b : 
  ( n1320 ) ? WR_XRAM_ADDR_0c : 
  ( n1315 ) ? WR_XRAM_ADDR_0d : 
  ( n1323 ) ? WR_XRAM_ADDR_0e : 
  ( n1325 ) ? WR_XRAM_ADDR_0f : 
  ( WR_XRAM_ADDR );
assign WR_XRAM_EN_next = 
  ( n1316 ) ? WR_XRAM_EN_00 : 
  ( n1313 ) ? WR_XRAM_EN_01 : 
  ( n1317 ) ? WR_XRAM_EN_02 : 
  ( n1318 ) ? WR_XRAM_EN_03 : 
  ( n1309 ) ? WR_XRAM_EN_04 : 
  ( n1310 ) ? WR_XRAM_EN_05 : 
  ( n1311 ) ? WR_XRAM_EN_06 : 
  ( n1312 ) ? WR_XRAM_EN_07 : 
  ( n1319 ) ? WR_XRAM_EN_08 : 
  ( n1314 ) ? WR_XRAM_EN_09 : 
  ( n1321 ) ? WR_XRAM_EN_0a : 
  ( n1322 ) ? WR_XRAM_EN_0b : 
  ( n1320 ) ? WR_XRAM_EN_0c : 
  ( n1315 ) ? WR_XRAM_EN_0d : 
  ( n1323 ) ? WR_XRAM_EN_0e : 
  ( n1325 ) ? WR_XRAM_EN_0f : 
  ( WR_XRAM_EN );
assign aes_state_next = 
  ( n1316 ) ? aes_state_00 : 
  ( n1313 ) ? aes_state_01 : 
  ( n1317 ) ? aes_state_02 : 
  ( n1318 ) ? aes_state_03 : 
  ( n1309 ) ? aes_state_04 : 
  ( n1310 ) ? aes_state_05 : 
  ( n1311 ) ? aes_state_06 : 
  ( n1312 ) ? aes_state_07 : 
  ( n1319 ) ? aes_state_08 : 
  ( n1314 ) ? aes_state_09 : 
  ( n1321 ) ? aes_state_0a : 
  ( n1322 ) ? aes_state_0b : 
  ( n1320 ) ? aes_state_0c : 
  ( n1315 ) ? aes_state_0d : 
  ( n1323 ) ? aes_state_0e : 
  ( n1325 ) ? aes_state_0f : 
  ( aes_state );
assign aes_enc_data_next = 
  ( n1317 ) ? aes_enc_data_02 : 
  ( n1311 ) ? aes_enc_data_06 : 
  ( n1321 ) ? aes_enc_data_0a : 
  ( n1323 ) ? aes_enc_data_0e : 
  ( aes_enc_data );
assign sha_state_next = 
  ( n1316 ) ? sha_state_00 : 
  ( n1313 ) ? sha_state_01 : 
  ( n1317 ) ? sha_state_02 : 
  ( n1318 ) ? sha_state_03 : 
  ( n1309 ) ? sha_state_04 : 
  ( n1310 ) ? sha_state_05 : 
  ( n1311 ) ? sha_state_06 : 
  ( n1312 ) ? sha_state_07 : 
  ( n1319 ) ? sha_state_08 : 
  ( n1314 ) ? sha_state_09 : 
  ( n1321 ) ? sha_state_0a : 
  ( n1322 ) ? sha_state_0b : 
  ( n1320 ) ? sha_state_0c : 
  ( n1315 ) ? sha_state_0d : 
  ( n1323 ) ? sha_state_0e : 
  ( n1325 ) ? sha_state_0f : 
  ( sha_state );
assign sha_digest_next = 
  ( n1316 ) ? sha_digest_00 : 
  ( n1313 ) ? sha_digest_01 : 
  ( n1317 ) ? sha_digest_02 : 
  ( n1318 ) ? sha_digest_03 : 
  ( n1309 ) ? sha_digest_04 : 
  ( n1310 ) ? sha_digest_05 : 
  ( n1311 ) ? sha_digest_06 : 
  ( n1312 ) ? sha_digest_07 : 
  ( n1319 ) ? sha_digest_08 : 
  ( n1314 ) ? sha_digest_09 : 
  ( n1321 ) ? sha_digest_0a : 
  ( n1322 ) ? sha_digest_0b : 
  ( n1320 ) ? sha_digest_0c : 
  ( n1315 ) ? sha_digest_0d : 
  ( n1323 ) ? sha_digest_0e : 
  ( n1325 ) ? sha_digest_0f : 
  ( sha_digest );

always @(posedge clk) begin
  if (rst) begin
    WR_XRAM_ADDR <= 16'h0;
    WR_XRAM_EN <= 0;
    aes_addr <= 16'h0;
    aes_bytes_processed <= 16'h0;
    aes_ctr <= 128'h0;
    aes_enc_data <= 128'h0;
    aes_key0 <= 128'h0;
    aes_key1 <= 128'h0;
    aes_len <= 16'h0;
    aes_read_data <= 128'h0;
    aes_state <= 8'h0;
    dataout <= 8'h0;
    sha_bytes_processed <= 16'h0;
    sha_digest <= 160'h0;
    sha_len <= 16'h0;
    sha_rdaddr <= 16'h0;
    sha_read_data <= 512'h0;
    sha_state <= 8'h0;
    sha_wraddr <= 16'h0;
  end
  else begin
    if (step) begin
      sha_read_data <= sha_read_data_next;
      aes_read_data <= aes_read_data_next;
      sha_rdaddr <= sha_rdaddr_next;
      aes_addr <= aes_addr_next;
      aes_ctr <= aes_ctr_next;
      aes_bytes_processed <= aes_bytes_processed_next;
      sha_len <= sha_len_next;
      aes_key1 <= aes_key1_next;
      aes_key0 <= aes_key0_next;
      aes_len <= aes_len_next;
      sha_bytes_processed <= sha_bytes_processed_next;
      sha_wraddr <= sha_wraddr_next;
      dataout <= dataout_next;
      WR_XRAM_ADDR <= WR_XRAM_ADDR_next;
      WR_XRAM_EN <= WR_XRAM_EN_next;
      aes_state <= aes_state_next;
      aes_enc_data <= aes_enc_data_next;
      sha_state <= sha_state_next;
      sha_digest <= sha_digest_next;
    end
  end
end

endmodule
