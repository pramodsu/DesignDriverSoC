module oc8051_xiommu_tb();

reg clk, rst;

reg proc_wr = 0, proc_stb = 0;
reg [7:0] proc_data_in = 0;
reg [15:0] proc_addr = 0;

reg [63:0] input_sha_func_0 = 0;
reg [63:0] input_sha_func_1 = 0;
reg [31:0] input_sha_func_2 = 0;
reg [63:0] input_sha_func_3 = 0;
reg [63:0] input_sha_func_4 = 0;
reg [31:0] input_sha_func_5 = 0;
reg [63:0] input_aes_func_6 = 0;
reg [63:0] input_aes_func_7 = 0;
reg [63:0] input_sha_func_8 = 0;
reg [63:0] input_sha_func_9 = 0;
reg [31:0] input_sha_func_10 = 0;
reg [63:0] input_sha_func_11 = 0;
reg [63:0] input_sha_func_12 = 0;
reg [31:0] input_sha_func_13 = 0;
reg [63:0] input_sha_func_14 = 0;
reg [63:0] input_sha_func_15 = 0;
reg [31:0] input_sha_func_16 = 0;
reg [63:0] input_sha_func_17 = 0;
reg [63:0] input_sha_func_18 = 0;
reg [31:0] input_sha_func_19 = 0;
reg [63:0] input_sha_func_20 = 0;
reg [63:0] input_sha_func_21 = 0;
reg [31:0] input_sha_func_22 = 0;
reg [63:0] input_aes_func_23 = 0;
reg [63:0] input_aes_func_24 = 0;
reg [63:0] input_sha_func_25 = 0;
reg [63:0] input_sha_func_26 = 0;
reg [31:0] input_sha_func_27 = 0;
reg [63:0] input_sha_func_28 = 0;
reg [63:0] input_sha_func_29 = 0;
reg [31:0] input_sha_func_30 = 0;
reg [63:0] input_sha_func_31 = 0;
reg [63:0] input_sha_func_32 = 0;
reg [31:0] input_sha_func_33 = 0;
reg [63:0] input_sha_func_34 = 0;
reg [63:0] input_sha_func_35 = 0;
reg [31:0] input_sha_func_36 = 0;
reg [63:0] input_aes_func_37 = 0;
reg [63:0] input_aes_func_38 = 0;
reg [63:0] input_sha_func_39 = 0;
reg [63:0] input_sha_func_40 = 0;
reg [31:0] input_sha_func_41 = 0;
reg [63:0] input_sha_func_42 = 0;
reg [63:0] input_sha_func_43 = 0;
reg [31:0] input_sha_func_44 = 0;
reg [63:0] input_sha_func_45 = 0;
reg [63:0] input_sha_func_46 = 0;
reg [31:0] input_sha_func_47 = 0;
reg [63:0] input_sha_func_48 = 0;
reg [63:0] input_sha_func_49 = 0;
reg [31:0] input_sha_func_50 = 0;
reg [63:0] input_aes_func_51 = 0;
reg [63:0] input_aes_func_52 = 0;
reg [63:0] input_sha_func_53 = 0;
reg [63:0] input_sha_func_54 = 0;
reg [31:0] input_sha_func_55 = 0;

reg [7:0] RD_xram_0 = 0;
reg [7:0] RD_xram_1 = 0;
reg [7:0] RD_xram_2 = 0;
reg [7:0] RD_xram_3 = 0;
reg [7:0] RD_xram_4 = 0;
reg [7:0] RD_xram_5 = 0;
reg [7:0] RD_xram_6 = 0;
reg [7:0] RD_xram_7 = 0;
reg [7:0] RD_xram_8 = 0;
reg [7:0] RD_xram_9 = 0;
reg [7:0] RD_xram_10 = 0;
reg [7:0] RD_xram_11 = 0;
reg [7:0] RD_xram_12 = 0;
reg [7:0] RD_xram_13 = 0;
reg [7:0] RD_xram_14 = 0;
reg [7:0] RD_xram_15 = 0;
reg [7:0] RD_xram_16 = 0;
reg [7:0] RD_xram_17 = 0;
reg [7:0] RD_xram_18 = 0;
reg [7:0] RD_xram_19 = 0;
reg [7:0] RD_xram_20 = 0;
reg [7:0] RD_xram_21 = 0;
reg [7:0] RD_xram_22 = 0;
reg [7:0] RD_xram_23 = 0;
reg [7:0] RD_xram_24 = 0;
reg [7:0] RD_xram_25 = 0;
reg [7:0] RD_xram_26 = 0;
reg [7:0] RD_xram_27 = 0;
reg [7:0] RD_xram_28 = 0;
reg [7:0] RD_xram_29 = 0;
reg [7:0] RD_xram_30 = 0;
reg [7:0] RD_xram_31 = 0;
reg [7:0] RD_xram_32 = 0;
reg [7:0] RD_xram_33 = 0;
reg [7:0] RD_xram_34 = 0;
reg [7:0] RD_xram_35 = 0;
reg [7:0] RD_xram_36 = 0;
reg [7:0] RD_xram_37 = 0;
reg [7:0] RD_xram_38 = 0;
reg [7:0] RD_xram_39 = 0;
reg [7:0] RD_xram_40 = 0;
reg [7:0] RD_xram_41 = 0;
reg [7:0] RD_xram_42 = 0;
reg [7:0] RD_xram_43 = 0;
reg [7:0] RD_xram_44 = 0;
reg [7:0] RD_xram_45 = 0;
reg [7:0] RD_xram_46 = 0;
reg [7:0] RD_xram_47 = 0;
reg [7:0] RD_xram_48 = 0;
reg [7:0] RD_xram_49 = 0;
reg [7:0] RD_xram_50 = 0;
reg [7:0] RD_xram_51 = 0;
reg [7:0] RD_xram_52 = 0;
reg [7:0] RD_xram_53 = 0;
reg [7:0] RD_xram_54 = 0;
reg [7:0] RD_xram_55 = 0;
reg [7:0] RD_xram_56 = 0;
reg [7:0] RD_xram_57 = 0;
reg [7:0] RD_xram_58 = 0;
reg [7:0] RD_xram_59 = 0;
reg [7:0] RD_xram_60 = 0;
reg [7:0] RD_xram_61 = 0;
reg [7:0] RD_xram_62 = 0;
reg [7:0] RD_xram_63 = 0;
reg [7:0] RD_xram_64 = 0;
reg [7:0] RD_xram_65 = 0;
reg [7:0] RD_xram_66 = 0;
reg [7:0] RD_xram_67 = 0;
reg [7:0] RD_xram_68 = 0;
reg [7:0] RD_xram_69 = 0;
reg [7:0] RD_xram_70 = 0;
reg [7:0] RD_xram_71 = 0;
reg [7:0] RD_xram_72 = 0;
reg [7:0] RD_xram_73 = 0;
reg [7:0] RD_xram_74 = 0;
reg [7:0] RD_xram_75 = 0;
reg [7:0] RD_xram_76 = 0;
reg [7:0] RD_xram_77 = 0;
reg [7:0] RD_xram_78 = 0;
reg [7:0] RD_xram_79 = 0;
reg [7:0] RD_xram_80 = 0;

reg nondet_memwrite_choice_0 = 0;
reg nondet_memwrite_choice_1 = 0;
reg nondet_memwrite_choice_2 = 0;
reg nondet_memwrite_choice_3 = 0;
reg nondet_memwrite_choice_4 = 0;
reg nondet_memwrite_choice_5 = 0;
reg nondet_memwrite_choice_6 = 0;
reg nondet_memwrite_choice_7 = 0;
reg nondet_memwrite_choice_8 = 0;
reg nondet_memwrite_choice_9 = 0;
reg nondet_memwrite_choice_10 = 0;
reg nondet_memwrite_choice_11 = 0;
reg nondet_memwrite_choice_12 = 0;
reg nondet_memwrite_choice_13 = 0;
reg nondet_memwrite_choice_14 = 0;
reg nondet_memwrite_choice_15 = 0;
reg nondet_memwrite_choice_16 = 0;
reg nondet_memwrite_choice_17 = 0;
reg nondet_memwrite_choice_18 = 0;
reg nondet_memwrite_choice_19 = 0;
reg nondet_memwrite_choice_20 = 0;
reg nondet_memwrite_choice_21 = 0;
reg nondet_memwrite_choice_22 = 0;
reg nondet_memwrite_choice_23 = 0;
reg nondet_memwrite_choice_24 = 0;
reg nondet_memwrite_choice_25 = 0;
reg nondet_memwrite_choice_26 = 0;
reg nondet_memwrite_choice_27 = 0;
reg nondet_memwrite_choice_28 = 0;
reg nondet_memwrite_choice_29 = 0;
reg nondet_memwrite_choice_30 = 0;
reg nondet_memwrite_choice_31 = 0;
reg nondet_memwrite_choice_32 = 0;
reg nondet_memwrite_choice_33 = 0;
reg nondet_memwrite_choice_34 = 0;
reg nondet_memwrite_choice_35 = 0;
reg nondet_memwrite_choice_36 = 0;
reg nondet_memwrite_choice_37 = 0;
reg nondet_memwrite_choice_38 = 0;
reg nondet_memwrite_choice_39 = 0;
reg nondet_memwrite_choice_40 = 0;
reg nondet_memwrite_choice_41 = 0;
reg nondet_memwrite_choice_42 = 0;
reg nondet_memwrite_choice_43 = 0;
reg nondet_memwrite_choice_44 = 0;
reg nondet_memwrite_choice_45 = 0;
reg nondet_memwrite_choice_46 = 0;
reg nondet_memwrite_choice_47 = 0;
reg nondet_memwrite_choice_48 = 0;
reg nondet_memwrite_choice_49 = 0;
reg nondet_memwrite_choice_50 = 0;
reg nondet_memwrite_choice_51 = 0;
reg nondet_memwrite_choice_52 = 0;
reg nondet_memwrite_choice_53 = 0;
reg nondet_memwrite_choice_54 = 0;
reg nondet_memwrite_choice_55 = 0;
reg nondet_memwrite_choice_56 = 0;
reg nondet_memwrite_choice_57 = 0;
reg nondet_memwrite_choice_58 = 0;
reg nondet_memwrite_choice_59 = 0;
reg nondet_memwrite_choice_60 = 0;
reg nondet_memwrite_choice_61 = 0;
reg nondet_memwrite_choice_62 = 0;
reg nondet_memwrite_choice_63 = 0;
reg nondet_memwrite_choice_64 = 0;
reg nondet_memwrite_choice_65 = 0;
reg nondet_memwrite_choice_66 = 0;
reg nondet_memwrite_choice_67 = 0;
reg nondet_memwrite_choice_68 = 0;
reg nondet_memwrite_choice_69 = 0;
reg nondet_memwrite_choice_70 = 0;
reg nondet_memwrite_choice_71 = 0;
reg nondet_memwrite_choice_72 = 0;
reg nondet_memwrite_choice_73 = 0;
reg nondet_memwrite_choice_74 = 0;
reg nondet_memwrite_choice_75 = 0;
reg nondet_memwrite_choice_76 = 0;
reg nondet_memwrite_choice_77 = 0;
reg nondet_memwrite_choice_78 = 0;
reg nondet_memwrite_choice_79 = 0;
reg nondet_memwrite_choice_80 = 0;
reg nondet_memwrite_choice_81 = 0;
reg nondet_memwrite_choice_82 = 0;
reg nondet_memwrite_choice_83 = 0;
reg nondet_memwrite_choice_84 = 0;
reg nondet_memwrite_choice_85 = 0;
reg nondet_memwrite_choice_86 = 0;
reg nondet_memwrite_choice_87 = 0;
reg nondet_memwrite_choice_88 = 0;
reg nondet_memwrite_choice_89 = 0;
reg nondet_memwrite_choice_90 = 0;
reg nondet_memwrite_choice_91 = 0;
reg nondet_memwrite_choice_92 = 0;
reg nondet_memwrite_choice_93 = 0;
reg nondet_memwrite_choice_94 = 0;
reg nondet_memwrite_choice_95 = 0;
reg nondet_memwrite_choice_96 = 0;
reg nondet_memwrite_choice_97 = 0;
reg nondet_memwrite_choice_98 = 0;
reg nondet_memwrite_choice_99 = 0;
reg nondet_memwrite_choice_100 = 0;
reg nondet_memwrite_choice_101 = 0;
reg nondet_memwrite_choice_102 = 0;
reg nondet_memwrite_choice_103 = 0;
reg nondet_memwrite_choice_104 = 0;
reg nondet_memwrite_choice_105 = 0;
reg nondet_memwrite_choice_106 = 0;
reg nondet_memwrite_choice_107 = 0;
reg nondet_memwrite_choice_108 = 0;
reg nondet_memwrite_choice_109 = 0;
reg nondet_memwrite_choice_110 = 0;
reg nondet_memwrite_choice_111 = 0;
reg nondet_memwrite_choice_112 = 0;
reg nondet_memwrite_choice_113 = 0;
reg nondet_memwrite_choice_114 = 0;
reg nondet_memwrite_choice_115 = 0;
reg nondet_memwrite_choice_116 = 0;
reg nondet_memwrite_choice_117 = 0;
reg nondet_memwrite_choice_118 = 0;
reg nondet_memwrite_choice_119 = 0;

wire property_invalid_aes_state;
wire property_invalid_sha_state;


initial
begin
  clk = 1;
  forever #100 clk <= ~clk;
end

initial
begin
  $dumpfile("run2.vcd");
  $dumpvars(0,oc8051_xiommu_tb);
  rst = 1'b1;
  #2001;
  rst = 1'b0;

`include "xiommu_cex.v"

  #80000
  $display("time ",$time, "; end of time\n");
  $finish;
end

oc8051_xiommu_gm_top oc8051_xiommu_gm_top_i(
    .clk(clk),
    .rst(rst),
    .proc_wr(proc_wr), 
    .proc_stb(proc_stb),
    .proc_addr(proc_addr), 
    .proc_data_in(proc_data_in), 

    .input_sha_func_0(input_sha_func_0), .input_sha_func_1(input_sha_func_1), .input_sha_func_2(input_sha_func_2), .input_sha_func_3(input_sha_func_3), .input_sha_func_4(input_sha_func_4),
    .input_sha_func_5(input_sha_func_5), .input_aes_func_6(input_aes_func_6), .input_aes_func_7(input_aes_func_7), .input_sha_func_8(input_sha_func_8), .input_sha_func_9(input_sha_func_9),
    .input_sha_func_10(input_sha_func_10), .input_sha_func_11(input_sha_func_11), .input_sha_func_12(input_sha_func_12), .input_sha_func_13(input_sha_func_13), .input_sha_func_14(input_sha_func_14),
    .input_sha_func_15(input_sha_func_15), .input_sha_func_16(input_sha_func_16), .input_sha_func_17(input_sha_func_17), .input_sha_func_18(input_sha_func_18), .input_sha_func_19(input_sha_func_19),
    .input_sha_func_20(input_sha_func_20), .input_sha_func_21(input_sha_func_21), .input_sha_func_22(input_sha_func_22), .input_aes_func_23(input_aes_func_23), .input_aes_func_24(input_aes_func_24),
    .input_sha_func_25(input_sha_func_25), .input_sha_func_26(input_sha_func_26), .input_sha_func_27(input_sha_func_27), .input_sha_func_28(input_sha_func_28), .input_sha_func_29(input_sha_func_29),
    .input_sha_func_30(input_sha_func_30), .input_sha_func_31(input_sha_func_31), .input_sha_func_32(input_sha_func_32), .input_sha_func_33(input_sha_func_33), .input_sha_func_34(input_sha_func_34),
    .input_sha_func_35(input_sha_func_35), .input_sha_func_36(input_sha_func_36), .input_aes_func_37(input_aes_func_37), .input_aes_func_38(input_aes_func_38), .input_sha_func_39(input_sha_func_39),
    .input_sha_func_40(input_sha_func_40), .input_sha_func_41(input_sha_func_41), .input_sha_func_42(input_sha_func_42), .input_sha_func_43(input_sha_func_43), .input_sha_func_44(input_sha_func_44),
    .input_sha_func_45(input_sha_func_45), .input_sha_func_46(input_sha_func_46), .input_sha_func_47(input_sha_func_47), .input_sha_func_48(input_sha_func_48), .input_sha_func_49(input_sha_func_49),
    .input_sha_func_50(input_sha_func_50), .input_aes_func_51(input_aes_func_51), .input_aes_func_52(input_aes_func_52), .input_sha_func_53(input_sha_func_53), .input_sha_func_54(input_sha_func_54),
    .input_sha_func_55(input_sha_func_55),

    .RD_xram_0(RD_xram_0), .RD_xram_1(RD_xram_1), .RD_xram_2(RD_xram_2),
    .RD_xram_3(RD_xram_3), .RD_xram_4(RD_xram_4), .RD_xram_5(RD_xram_5),
    .RD_xram_6(RD_xram_6), .RD_xram_7(RD_xram_7), .RD_xram_8(RD_xram_8),
    .RD_xram_9(RD_xram_9), .RD_xram_10(RD_xram_10), .RD_xram_11(RD_xram_11),
    .RD_xram_12(RD_xram_12), .RD_xram_13(RD_xram_13), .RD_xram_14(RD_xram_14),
    .RD_xram_15(RD_xram_15), .RD_xram_16(RD_xram_16), .RD_xram_17(RD_xram_17),
    .RD_xram_18(RD_xram_18), .RD_xram_19(RD_xram_19), .RD_xram_20(RD_xram_20),
    .RD_xram_21(RD_xram_21), .RD_xram_22(RD_xram_22), .RD_xram_23(RD_xram_23),
    .RD_xram_24(RD_xram_24), .RD_xram_25(RD_xram_25), .RD_xram_26(RD_xram_26),
    .RD_xram_27(RD_xram_27), .RD_xram_28(RD_xram_28), .RD_xram_29(RD_xram_29),
    .RD_xram_30(RD_xram_30), .RD_xram_31(RD_xram_31), .RD_xram_32(RD_xram_32),
    .RD_xram_33(RD_xram_33), .RD_xram_34(RD_xram_34), .RD_xram_35(RD_xram_35),
    .RD_xram_36(RD_xram_36), .RD_xram_37(RD_xram_37), .RD_xram_38(RD_xram_38),
    .RD_xram_39(RD_xram_39), .RD_xram_40(RD_xram_40), .RD_xram_41(RD_xram_41),
    .RD_xram_42(RD_xram_42), .RD_xram_43(RD_xram_43), .RD_xram_44(RD_xram_44),
    .RD_xram_45(RD_xram_45), .RD_xram_46(RD_xram_46), .RD_xram_47(RD_xram_47),
    .RD_xram_48(RD_xram_48), .RD_xram_49(RD_xram_49), .RD_xram_50(RD_xram_50),
    .RD_xram_51(RD_xram_51), .RD_xram_52(RD_xram_52), .RD_xram_53(RD_xram_53),
    .RD_xram_54(RD_xram_54), .RD_xram_55(RD_xram_55), .RD_xram_56(RD_xram_56),
    .RD_xram_57(RD_xram_57), .RD_xram_58(RD_xram_58), .RD_xram_59(RD_xram_59),
    .RD_xram_60(RD_xram_60), .RD_xram_61(RD_xram_61), .RD_xram_62(RD_xram_62),
    .RD_xram_63(RD_xram_63), .RD_xram_64(RD_xram_64), .RD_xram_65(RD_xram_65),
    .RD_xram_66(RD_xram_66), .RD_xram_67(RD_xram_67), .RD_xram_68(RD_xram_68),
    .RD_xram_69(RD_xram_69), .RD_xram_70(RD_xram_70), .RD_xram_71(RD_xram_71),
    .RD_xram_72(RD_xram_72), .RD_xram_73(RD_xram_73), .RD_xram_74(RD_xram_74),
    .RD_xram_75(RD_xram_75), .RD_xram_76(RD_xram_76), .RD_xram_77(RD_xram_77),
    .RD_xram_78(RD_xram_78), .RD_xram_79(RD_xram_79), .RD_xram_80(RD_xram_80),

    .nondet_memwrite_choice_0(nondet_memwrite_choice_0),
    .nondet_memwrite_choice_1(nondet_memwrite_choice_1),
    .nondet_memwrite_choice_2(nondet_memwrite_choice_2),
    .nondet_memwrite_choice_3(nondet_memwrite_choice_3),
    .nondet_memwrite_choice_4(nondet_memwrite_choice_4),
    .nondet_memwrite_choice_5(nondet_memwrite_choice_5),
    .nondet_memwrite_choice_6(nondet_memwrite_choice_6),
    .nondet_memwrite_choice_7(nondet_memwrite_choice_7),
    .nondet_memwrite_choice_8(nondet_memwrite_choice_8),
    .nondet_memwrite_choice_9(nondet_memwrite_choice_9),
    .nondet_memwrite_choice_10(nondet_memwrite_choice_10),
    .nondet_memwrite_choice_11(nondet_memwrite_choice_11),
    .nondet_memwrite_choice_12(nondet_memwrite_choice_12),
    .nondet_memwrite_choice_13(nondet_memwrite_choice_13),
    .nondet_memwrite_choice_14(nondet_memwrite_choice_14),
    .nondet_memwrite_choice_15(nondet_memwrite_choice_15),
    .nondet_memwrite_choice_16(nondet_memwrite_choice_16),
    .nondet_memwrite_choice_17(nondet_memwrite_choice_17),
    .nondet_memwrite_choice_18(nondet_memwrite_choice_18),
    .nondet_memwrite_choice_19(nondet_memwrite_choice_19),
    .nondet_memwrite_choice_20(nondet_memwrite_choice_20),
    .nondet_memwrite_choice_21(nondet_memwrite_choice_21),
    .nondet_memwrite_choice_22(nondet_memwrite_choice_22),
    .nondet_memwrite_choice_23(nondet_memwrite_choice_23),
    .nondet_memwrite_choice_24(nondet_memwrite_choice_24),
    .nondet_memwrite_choice_25(nondet_memwrite_choice_25),
    .nondet_memwrite_choice_26(nondet_memwrite_choice_26),
    .nondet_memwrite_choice_27(nondet_memwrite_choice_27),
    .nondet_memwrite_choice_28(nondet_memwrite_choice_28),
    .nondet_memwrite_choice_29(nondet_memwrite_choice_29),
    .nondet_memwrite_choice_30(nondet_memwrite_choice_30),
    .nondet_memwrite_choice_31(nondet_memwrite_choice_31),
    .nondet_memwrite_choice_32(nondet_memwrite_choice_32),
    .nondet_memwrite_choice_33(nondet_memwrite_choice_33),
    .nondet_memwrite_choice_34(nondet_memwrite_choice_34),
    .nondet_memwrite_choice_35(nondet_memwrite_choice_35),
    .nondet_memwrite_choice_36(nondet_memwrite_choice_36),
    .nondet_memwrite_choice_37(nondet_memwrite_choice_37),
    .nondet_memwrite_choice_38(nondet_memwrite_choice_38),
    .nondet_memwrite_choice_39(nondet_memwrite_choice_39),
    .nondet_memwrite_choice_40(nondet_memwrite_choice_40),
    .nondet_memwrite_choice_41(nondet_memwrite_choice_41),
    .nondet_memwrite_choice_42(nondet_memwrite_choice_42),
    .nondet_memwrite_choice_43(nondet_memwrite_choice_43),
    .nondet_memwrite_choice_44(nondet_memwrite_choice_44),
    .nondet_memwrite_choice_45(nondet_memwrite_choice_45),
    .nondet_memwrite_choice_46(nondet_memwrite_choice_46),
    .nondet_memwrite_choice_47(nondet_memwrite_choice_47),
    .nondet_memwrite_choice_48(nondet_memwrite_choice_48),
    .nondet_memwrite_choice_49(nondet_memwrite_choice_49),
    .nondet_memwrite_choice_50(nondet_memwrite_choice_50),
    .nondet_memwrite_choice_51(nondet_memwrite_choice_51),
    .nondet_memwrite_choice_52(nondet_memwrite_choice_52),
    .nondet_memwrite_choice_53(nondet_memwrite_choice_53),
    .nondet_memwrite_choice_54(nondet_memwrite_choice_54),
    .nondet_memwrite_choice_55(nondet_memwrite_choice_55),
    .nondet_memwrite_choice_56(nondet_memwrite_choice_56),
    .nondet_memwrite_choice_57(nondet_memwrite_choice_57),
    .nondet_memwrite_choice_58(nondet_memwrite_choice_58),
    .nondet_memwrite_choice_59(nondet_memwrite_choice_59),
    .nondet_memwrite_choice_60(nondet_memwrite_choice_60),
    .nondet_memwrite_choice_61(nondet_memwrite_choice_61),
    .nondet_memwrite_choice_62(nondet_memwrite_choice_62),
    .nondet_memwrite_choice_63(nondet_memwrite_choice_63),
    .nondet_memwrite_choice_64(nondet_memwrite_choice_64),
    .nondet_memwrite_choice_65(nondet_memwrite_choice_65),
    .nondet_memwrite_choice_66(nondet_memwrite_choice_66),
    .nondet_memwrite_choice_67(nondet_memwrite_choice_67),
    .nondet_memwrite_choice_68(nondet_memwrite_choice_68),
    .nondet_memwrite_choice_69(nondet_memwrite_choice_69),
    .nondet_memwrite_choice_70(nondet_memwrite_choice_70),
    .nondet_memwrite_choice_71(nondet_memwrite_choice_71),
    .nondet_memwrite_choice_72(nondet_memwrite_choice_72),
    .nondet_memwrite_choice_73(nondet_memwrite_choice_73),
    .nondet_memwrite_choice_74(nondet_memwrite_choice_74),
    .nondet_memwrite_choice_75(nondet_memwrite_choice_75),
    .nondet_memwrite_choice_76(nondet_memwrite_choice_76),
    .nondet_memwrite_choice_77(nondet_memwrite_choice_77),
    .nondet_memwrite_choice_78(nondet_memwrite_choice_78),
    .nondet_memwrite_choice_79(nondet_memwrite_choice_79),
    .nondet_memwrite_choice_80(nondet_memwrite_choice_80),
    .nondet_memwrite_choice_81(nondet_memwrite_choice_81),
    .nondet_memwrite_choice_82(nondet_memwrite_choice_82),
    .nondet_memwrite_choice_83(nondet_memwrite_choice_83),
    .nondet_memwrite_choice_84(nondet_memwrite_choice_84),
    .nondet_memwrite_choice_85(nondet_memwrite_choice_85),
    .nondet_memwrite_choice_86(nondet_memwrite_choice_86),
    .nondet_memwrite_choice_87(nondet_memwrite_choice_87),
    .nondet_memwrite_choice_88(nondet_memwrite_choice_88),
    .nondet_memwrite_choice_89(nondet_memwrite_choice_89),
    .nondet_memwrite_choice_90(nondet_memwrite_choice_90),
    .nondet_memwrite_choice_91(nondet_memwrite_choice_91),
    .nondet_memwrite_choice_92(nondet_memwrite_choice_92),
    .nondet_memwrite_choice_93(nondet_memwrite_choice_93),
    .nondet_memwrite_choice_94(nondet_memwrite_choice_94),
    .nondet_memwrite_choice_95(nondet_memwrite_choice_95),
    .nondet_memwrite_choice_96(nondet_memwrite_choice_96),
    .nondet_memwrite_choice_97(nondet_memwrite_choice_97),
    .nondet_memwrite_choice_98(nondet_memwrite_choice_98),
    .nondet_memwrite_choice_99(nondet_memwrite_choice_99),
    .nondet_memwrite_choice_100(nondet_memwrite_choice_100),
    .nondet_memwrite_choice_101(nondet_memwrite_choice_101),
    .nondet_memwrite_choice_102(nondet_memwrite_choice_102),
    .nondet_memwrite_choice_103(nondet_memwrite_choice_103),
    .nondet_memwrite_choice_104(nondet_memwrite_choice_104),
    .nondet_memwrite_choice_105(nondet_memwrite_choice_105),
    .nondet_memwrite_choice_106(nondet_memwrite_choice_106),
    .nondet_memwrite_choice_107(nondet_memwrite_choice_107),
    .nondet_memwrite_choice_108(nondet_memwrite_choice_108),
    .nondet_memwrite_choice_109(nondet_memwrite_choice_109),
    .nondet_memwrite_choice_110(nondet_memwrite_choice_110),
    .nondet_memwrite_choice_111(nondet_memwrite_choice_111),
    .nondet_memwrite_choice_112(nondet_memwrite_choice_112),
    .nondet_memwrite_choice_113(nondet_memwrite_choice_113),
    .nondet_memwrite_choice_114(nondet_memwrite_choice_114),
    .nondet_memwrite_choice_115(nondet_memwrite_choice_115),
    .nondet_memwrite_choice_116(nondet_memwrite_choice_116),
    .nondet_memwrite_choice_117(nondet_memwrite_choice_117),
    .nondet_memwrite_choice_118(nondet_memwrite_choice_118),
    .nondet_memwrite_choice_119(nondet_memwrite_choice_119),

    .property_invalid_aes_state(property_invalid_aes_state),
    .property_invalid_sha_state(property_invalid_sha_state)
);

endmodule
